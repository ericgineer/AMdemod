`timescale 1ns/1ns

`define width 72

module CIC(
	input wire               clk,
	input wire               rst,
	input wire        [15:0] decimation_ratio,
	input wire signed [7:0]  d_in,
	output reg signed [7:0]  d_out,
	output reg 				 d_clk
);

reg signed [`width-1:0] d_tmp, d_d_tmp;


// Integrator stage registers

reg signed [`width-1:0]  d1, d_d1;
reg signed [`width-1:0]  d2, d_d2;
reg signed [`width-1:0] d3, d_d3;
reg signed [`width-1:0] d4, d_d4;
reg signed [`width-1:0] d5, d_d5;

// Comb stage registers

reg signed [`width-1:0] d6, d_d6;
reg signed [`width-1:0] d7, d_d7;
reg signed [`width-1:0] d8, d_d8;
reg signed [`width-1:0] d9, d_d9;
reg signed [`width-1:0] d10;

reg [15:0] count;

 
	always @(posedge clk)
	begin
		if (rst)
		begin
			d1 <= 0;
			d2 <= 0;
			d3 <= 0;
			d4 <= 0;
			d5 <= 0;
			d6 <= 0;
			d7 <= 0;
			d8 <= 0;
			d9 <= 0;
			d10 <= 0;
			d_out <= 0;
			
			d_d1 <= 0;
			d_d2 <= 0;
			d_d3 <= 0;
			d_d4 <= 0;
			d_d5 <= 0;
			d_d6 <= 0;
			d_d7 <= 0;
			d_d8 <= 0;
			d_d9 <= 0;
			count <= 0;
			d_clk <= 1'b0;
		end else
		begin
			// Integrator section
			d1 <= d_in + d_d1;
			d_d1 <= d1;
			
			d2 <= d1 + d_d2;
			d_d2 <= d2;
			
			d3 <= d2 + d_d3;
			d_d3 <= d3;
			
			d4 <= d3 + d_d4;
			d_d4 <= d4;
			
			d5 <= d4 + d_d5;
			d_d5 <= d5;
			
			// Decimation
			
			if (count == decimation_ratio - 1)
			begin
				count <= 16'b0;
				d_tmp <= d5;
				d_clk <= 1'b1;
			end else if (count == decimation_ratio >> 1)
			begin
				d_clk <= 1'b0;
				count <= count + 1;
			end else
				count <= count + 1;
		end
	end
	
	always @(posedge d_clk)  // Comb section running at output rate
	begin	
		// Comb section
		d_d_tmp <= d_tmp;
		
		d6 <= d_tmp - d_d_tmp;
		d_d6 <= d6;

		d7 <= d6 - d_d6;
		d_d7 <= d7;

		d8 <= d7 - d_d7;
		d_d8 <= d8;

		d9 <= d8 - d_d8;
		d_d9 <= d9;

		d10 <= d9 - d_d9;
		
		d_out <= d10 >>> (`width - 8);
	end								
endmodule
