��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I���t譈ȟ�R���ZK���/�%�G�%�^5�[0σ20#�>�|2T�p�}���~�B��6%H�&�\*�j�K�Fr$H{=Ǆ/�MbO����PLH��#S�0rȚ����r�/{�H�+������V��*� �w����� �	��$�J�v^|�	�tOk((�)�ɩ÷�3M��%v#�R�1�oJt���d�b2�{�(Al��b��������N]���kŤ�`cB���!q"2�m=:�Ұ��q��EK$:��\�E����z���<��3l2j��a�7]P��MD�a��Z0ɖ�ԇ�V�?�tU��`�'���sr5�.�TxJ�_\Iܳ�Y���)�$�}�6�#���Hh�^毪\���a�h�a@��#ń�����υj8hE�h����O��{A����,6���2�
 ���Aʠ����!ɨ�O{�a�<�˨�VB��*0`P�G�ʭ�&�z6���ytcE�k�1�RzЯ��jh#֦��Gp��c�q�Z����h�H81<��.i�C��/���Rc悴�F㙆:�)Z(cΘ�V� ��"��?�{�&j���b��
� PVMX���L6�5������?�C�0M��Bv�:ˬ+���X;�������ů��F�,Å�5���M�K��nVAh�04��;,�p5�g��C�v�V��p�/�q� ��#��8T�0*�*�:M���_Ϥ|���nAZ� ��:��D�*��V ��"��a~�x�(�^,�{�P&�FY���-nY���sw7��[�('/+�TV�����x��u�/I!�����4�u><*����{��;�/Т~����[��qs݉^<л� y�,�8�B	3�UC�p���IT�%�ڗ���/e�>�$����>��/k�bZ p��h�
��5{�8-`��ٌ�O�6����Wü ~Id�=\�a�����NZ���~8�>�c��BX��Ȭ�x�����̮#�-�]£(6P�	���x�zc�4AQ�J��c5�釻��v���^e0}��3���L��TH�����w&�s�f_���N2_�[��f�@�%З���_Z��g����PK����!��׫��,R��2vOY��EF�yDs1Q�1R)����o����Ds�7���x�<{��.f7j�!�q��B��/d�9rgW��h���%��F��ք[y�����\�b��C9ݽpW���j|O�Z��������(\(������:��)IH�&;>E����#�MxMC�.��r�%��L'ҧºCL�p)�¥�!��ؒg�Ӊ�����"������I\w���,�#V�����ֱ�������%�S8�I�M��ψ��De�,H�/�g9$��x��Dw�|��`K@~�)�uz��:ٞ�	��^�f�� t�#N"�?9k�0A9#�'����z��B�ٚ#8a��2�_IM潣��T8X�yK~��~l�Q����R�_CXj�t������7�K�em�(�n�`��\�g�6��1���c�Ǚ��S!k�Nx��J��PD�}���ߑ��c�����ի��.�mg��B박2璹e� E6A�l�R�Ma/6'���=��	E`�N]��T�s�ݦ��h<�˄R����_�.�����9G�$���N{�-t�.�)����JX\�]��$!�Eez�����IL�Ь����P�ʠu�T<~*��t\�:��o�ΩDؿ�`x&}h0�{]Q�x�rW���;��4��|K\�d� �U�?�0����Uj���p����f�p�~���U�]��V��}��o$�ֳ�L'���}m�{,����T��{G�G\t��3%�*b����A_��[Dk�f%��XD�Xy���m��k��NO���)���'�œ��B'��u�)�fT5�T&t\s_Qi���z;�/3T���U��5`߂�5�P�n7���S
@yY8Vn=���9Βt���7ӵ(,�-�Z��ΐ�gv�Ka,sիt\�1�g�M�U���A��]�� I� NWN�OZ�Eo{��H�T���(�X'�A�Q���8=As��z��{���Q
X�; ;c!�N�oI��xP��#�k���	�UP'iAD���]���m��F	��ܿ8A�>������M��k2��/�m6�F�Ƙ�o��B���3|�69���������������<V�Ǚ�H����+�J����[��nG6�=L)�zg����i @J!��~�]��&Y�I�C����Kt�D��L�6���oq2��ٶ2�q.c����]�UkX�y�<;u�ϧ(��|�5[!�"��C�A�9D��{Y�:^�`�R�k�����AQT���F�tOe`�}o���5|Ժ�d-h�x�+��?�G82jE���x�:�}� i�0K�D ���KU@�!P9]{�0>�G�Ҹ�X�[��/B��}��v�Ir�i	��șH�Ǻ5�a�]�v!��'TbW��w�=���Vl�v�C��^��Q�q���'<r�����Pu���a�j��
+�˞w�;E��{R'$���f*�y���0�a���(�/28^��hi��t�Eo�� X{�?����L�$V��ꮣ�0������!	��-�����ِ����26��S�W�~;�<�e�0��Et2�\��Vz���"��8�I~*Ahr���^XBFSi�$s�>���8RB�$�{w��t��X�g۸[c<Jɡ��Sz?d���4�%�f�i�F��$�sȧ�,~hEj.��b� �Nr�0πG$��C	�I�'�OGQ��2�JG{��@l?d&�[kH���3e��w�YM���!�dh�/h䥩<�p��0�t=1g̾�/1.r�����,��ż�YJ˭�<�|���x&�Rq��P�{�7���@~*0$;�M