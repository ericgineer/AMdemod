��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�����g��y�(.��H�^���z=ͦj�P@���I��_]�E�����U��@�iKAUu��z��}Kk�4�m�dC_�0w+�͹.a(:��D����ɿvw��s��=��PS?�8�\р��9ꌭ���:`��E=��8u3 ��;��\������k�@s���|������)���J �ꨣ�҇�6Q�?����G�����d�@hc͌o_� U���"U�4��ͯ�>���l?f�7h��z�U�]�\in�+4��l
[�W�*�鉪G��Nj�lzR�5�bV�����2���+�+�[��Q_#(�0h�9V�C��N���P����r��-���s�vw+�j����_	N���h��TY�j�N��x�8fy��_�OFZe3�e��CFY���@���$-9��wD��I�+�=�K���mI�>��D��>{NK�cM��e�Q����Tֵ�����H�)�|B��t��oXL��@��3�;F%�i���6�=���pKn�_�9^��3�fz[��_a���79��@b��n���,��{�M��EL��蒠�7Dr}u�bA�3m����{��Ȫ���4l�A��?v��(2N$���Sj[�=mm�?o��И#kg��2�~��Ui���X���dM⎷���4���`��`j`�A��xalC}C�?�Ło}�	ȭ�몽y��)x�ɏ��yx���9p]�\��DL+Xޙ��T_�d�=�C���)*9�A=;I"&d2`�Ȗ���8��t�F�.�ӆZe7�~*B!շX�UTc��O�!�熕j�h_��*L�K/�Һ���1��W���ٖx��ꐪV=LZ��(ҭG๑Z��e!x)�{>�n}��Ԓ�Z"0:������z7;�,I_K�Jl<��pkѨ�4k@@5Q�r�<�p�ZD
<Jc��=�*���.nH�,�!ws�ڲ�[�L��}�({r�+���y�|��P&���4B�VK�-�SE�A��K#��(P2l$!(��h����Ԥ�_�y08��h���y�e���H��Ũ�4����H@�떞_��d4�AY���zHB�fȋ�!�m�:�P�b���o
ȫ'q^E�	2tG���\ǡhi������ּ�!����!:]
.<1}2���6؀�	Xd����&D{��c�1E�RDY�W[ قs�c.)��M�ε��?;�pI�/�bە+}&��<Q�/MP}����ܥ�
)���M�{�s���j�A��-�c��ȸ���V�J`�f6cm��אD-�MՆ�[cL��/F�V/�b|�@���<pt\�F���,�f�Z}�~ߑ�.	����q������M��u]�@�"z᳢�m�ͥ�ҵ�YP4eY��z;��d���O85�4��+ne�H#�z���$���y8 Cu^�Ĵe�H�O,��"��V�Gٮ~F8��1S���h�����A(9x{Ӯ��� �=�?!���o~��8����2�/��X�y���+j��R/"�@\)M2���ɓ�t	;ɣ�]o��o�`��k��
@�~�	�P<N�e8��&t�t���� ��Լq	���RзޙE2׃�pP�a�?_L>�qڎ�CYu^1R��*�?�!��"5P��$hw����}�ܳZ�Ȧ�=�Sw��(4�����)0�©i:/���L����Ms��_��\"���lݽ�s�k��(�ES�u�
{��� �{��
�u�rx�;���,AlӀ�^�&P�G�S%>ba�.;0��WR\:�~��o��  <�-�V���
프 Y�&m��<Hy�	%�@9J��/��70�i�)o��U�}�}�17���Ql�|���E&ҬԨ4!�O�jm�,0��&��$5"d�\fEd�P��(wd�Lח6pUc���6�T�QM%�%C>�=����q>֛���L1!(��X���?n6{jc�z�"Uc�`\�=eG�T��W�����S�
I�]7��qei~z�����E�5�2*�"m�
�vT{�MM��E��V��A�hz�zU���U]nRB��RD����������L^Pi�����:��΍���wC
�iP˦�U;v�S5&� ��OA����`�z���ȷzJh���"��o�`�Β���^|n���,�Vy���.��_�1�?nC�N���ߛ ��fpNW�La9-�jBp|��H���B%T���ѽ�d���2�MRW��ꇗ�Ok	�AP���Vowx\�Reʅ�4�$пn�K��A9ҏ�5���$v�x�t����>��!�%�N�g��Ϳ�;�~�Ș|؏�5�Fg/��g���������l!f�ؾ���-���ۈ���XB�:�{o]/��d�6�q	c=~������go@����V��-����TCo6p�Jz��*J���Sj��nbZڛ���s{n�~A GX�%?wbe���r{GȬ���C/\%S}0g�@��½7"�O���XV��MI���%�6@��$
� ��|� ��4��mB�'�D�A��,�E�73<�|��+THh��Ę�vU�����^Uk������N�<K6$ߙ;��Q�����k�v�s{e���k*Gq��h�ߍ��RO�k���)�%1�l���T���{�6�j��0Vlճ?��O�������w�T�C���;/�h���(;�u���Z��O�(xCf>��JFA���Ǽ&�[����
Oh��O��m6��2�,��´1ߞ���f�\���R�3��l��~>�h}C���tAޘ�iO��b1�t�����pw��v�fp��Pt����Z�;\�6��߻.Z�S�8��@�]�{�-���Q�6�*�/�^�G�%�x'(GZ"����=X�OPJd@��7� �%(���dA���%����2�����K/�,��"F�"�4�����0	e;ɶ��ZDY������oΪ���������^e�]@v�7��3����Y���xTdC$�r�Ʊ�}�H���� ���T����۫�$u�� 3�afD�˲�������j��UB��
r`֬���f�敬��
�ć1�%�Qo5=)�^�d�U!|M�a�?�y��a�	���@�Ru.X)!ڷ����_ �.\�{�>�����&�L���}}��#b��˝�F�$R|�Zf͂��H��h��b�ڭx�ǖ�鍕��+�R��s��JQ(�5�Oh�`KNAv���lel�k�z�Y�����6�����s����]ܯ���P��K��8���#\"5�{
&oc�M�e�}%Ta��'0z�/	o�j�cj�I�UbH ��_L�G�[3�3�`����������2BȱĹ��ú�1���K�RqW��ޮ�UEP��kёT��xA�6LڟT���q7B�Y�PGB�\+�t�+�6�g���8.�}'�|5�g�#��y^^�?��������n�〒:џC����fM���q��ll�w�s.�&_'���9q���Բ����ޒ/ӑ�Ju��n�ϼ��-�*\e]���MJy��V9@��=�R���S�0�6��On�q��B �W̍e%aZkC�z�u��N�4���˄�#�"n��&O�<ho�Eh��b����i�#�Y,�3�g�H��XȪ'e`5N�H��� �k�'�o���+�Gv_ET]#����oѐ(m|'�Mo��p�&�$O�-�3�����{���ol+P����v�?���?Z�k>�-�F�u]��0WyM1}�N��BF�<��{� رd8��^o&���o^x�G?G:ʦ����°�1\2%`���]�O�O����*�� \� 9�3��y+���<�O�Z�wT[�Z���[ֿ;�5�UP�1�˨FOj����w���UP�MNJ���mO�$6c< C�K����X`���Լ�|�m��>������"��qٝ-J7H��E��+�h�RY���P������(��G r�$�@.4�~���RN��\N�1��1���W��M���y4|a�PER�M��}HJ�V\�Ov���Z+�I���I��"�����a&��,� �={|!]@YOk�T���^��@0�9^'�*�ɛ��w׃��u�M���
�%iP%�UY�i�q*�O�A"���Hx�<�ԍB��
�M��Z<j�H!��m+/�b�9�U�!څ	�I�f6��nn��m�I>�i۫� MT��M��� �^.��(��P�MϑgU�n�3#� �	F��u�X)�ǐ�7V�$Sd�s�$���cQ=�XC#�i��u� X±W�G���B|�]���1��k?,�`#����E�o,�ɣ���@~�u#o���D,�`)�$f�|$}}]>�{7e§�9K!T�4D	����>�o¬Z�
�[�<���������IѠ0ŕ��g ��46�h��VK�ڸ>�<B4�$ZB
'�Ty�Q�R�^��������3�����vn=4j5������ՌqβS���ok�'���,r��Pk밣)��N�%v��=si	�?�:�P-y��[`0\�����H_�1(���]Sfԃ״W%�(q'w�`ed�yQ��s㸰���z��zy��9�zV�@$��:�r*��+���h¨��� \�L���Y;+gǭq��♕l��A���ɂp/a\�@ho�d5���_���Fk�&���.�Vz�o����D,0������F���Cu�.x#u,�r���i�W.��^�KP�bB�θ2�Lf��C3"��`����r5�P#���,�U�΄%���~��G72�'�7<�פ^Y��7Jd֜�e�
��2ԞKb�o�D��|�C�ڗ�Rt©j"����m�]~ 萿B��Ouc>�-�����+���P����ɯ�G�{�%ٻ����l���"	qN�N�\�A�¾[������R�v_`$��[>���iXy����@�V�+z�p-�eN#u}D:�p����9~�H4�4G�ju��jT����8RY+�_6Y�NxU1Q	쏉w�۬��%l��=��B�Qe�챡\�=���] �7�d�g�L�9h5���06�ܠ�ox"%���)VP�UG�_��g�����ԨT!K»V���WM��"z�X|pLZ���P�n��^iC��3
�� �P�o�4�Z�1���$��< U((S�?Ȯ�ٍ��D�)ř�_��@}��V�xYX��|���_�As�Y{x���/��{�O�vh��Mh�$_�؇%�����[y�����Q(׌>oҴF��\uTVĨx�]��{��D&����dUR+�vA꠼�v �%�t�MK���}._��Ѽmkxb�42�%z�q��&��|6N��x�а!y]M3���6����R,�� �ST�_t7J�}����{�����^RԐr���O��V��F!}��ŗ��$ͥܕ�6�����=�3X����N�&1�"{&T���P�J�=<s��6�]�h#L�=5�<�㳄/˙��OP�#~��[;����)�A�x�����a��HP�+�wcѹ��>�=&�+�w�$j�p���g�?��D��7q�nn����xo���0Gy�؀wr��f��qAXʶ�mj�M`\z��U���'�c�!qٓ�� �2#�n/R�v���5-L� ໿=��Ÿ�n�G�1�OSќ���[��
8p�o��e��E؊��w	Q3.;1����	�7ٔD�!�9dd]����H��"QTM����	fڦ���C�T��Ư���a�s	��ð5����g>!9��bF�ܞ���;&?R+��-\�फ़�I�	��&������΂���C�x��,�X0�`�O�Dt7(r>?YzQ�/5qZӺ|Eچ��[��bf���nm^�Ȩ]X�eI� 6 Kt�uDh�JNS��{M�P�C`�@�@W���D�9�~��z���Re<[{�,-��x�)6���]Cp�x�q��x �,��Ӝ�2�A�Фe�{O�Hhlf��N��x+o�yX`0v�{}o��>*��z����Y��K+{����^p΄\(Z��^(�h�+�5�����R �jHÓ5U���~�r��W����z�],0>��e>y���S�#�pJ�)���ti��{Xw��#Y�X����kV�y3�}1�]J6B|�߷�I]�A�"x4[\ߚq=#���5��=±��j���K��5jy ~	�D��#e�[�B}��to(�^�1uk�����X�I~�����l�H�Ñ���kwY���=@jЯ�Qv�L$����j2?s�����nH��EP1���Q��~A˵���;<�����p��QM��C�#�sER�0�o�z})�nʯ��3������Xq����<y�WK?c7�o��$�t�T!*~�oJ��$�m�6�K��((�v��C�^�g���'��A�Cb�%?\5��y6J����
`3�T ��å����_l�@�[��9�� �CM���^�(�g��4��QD�b.�	���xNu:ɩ�
��aK^]�3�hU���<����A@[�;x��L�&B��( �Xg���o��Ԇ��A"�@��^[���_gP���3 �2Dx
��R-)�l���>��$&]���}m񆧹��gxN��OV�������8����~3��l��С�DO�Õ���g�(D�����Gtx��5�K������Z%�u:jk�xM�1�?/��~x��d�E�kP!��fyߡň�`_�F�BX����f�'ђ�Nu�o*LI$u��K�w�@6���ü{�~�rL/�ȹ��XXq��5�ȥY� �F��A_W&��B#��lǅ6!p��85�8�7��+�`S�.ʭޘ]6�X y_<o��1�|TJ6���c����y�}8 Y:������4��T)$|�����MgcG���L�mF_@���N��Cc�{0�
�lt�� y�Fk�}��UPXh�����'ʩ]WdZmo��蚃m��~�����[I��#�}q�j�[v�E<">�i�QL���;�@����gݻ������~;�)$��j�(~K�&8�[��{h]�%_P�߭�G��q#u��\���Q�{M����L�
���m�L@!��8%��J��g��8�A�\!�Pr n�9