��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��Mg9��X����6���
;gKd��Z{ferbwN�m��P5%�a9�/;�ۜlڿ�I0(��Z삥��*T;��3���*Hč�kOg��L.;v�ȫWr�_d!��H�0�/���d���Z$�OV���hà
�3���w�� ���;�	_�Ϲ�����\䌕+����0�l�HϿܠm?�Q��\�ՙ��o�Пoʻk����w�=P�=�C_��OF���S#v�8���#��J�|�H:�@�U[_��}^sK^���g��|�7��x/��_��N���1��6� 恲@�)�.� K�̟�҆H7�;8�w`����0P��8�G`5�Y|fd&Y����e�#B_�PxIkof>����y����뎒F@�}����������$ "$y*#�F����$4���ſ��Jqё�������ŶK��/��ʤ�����/�E�i^��L�AH��M���<�	��=�ր�_N�d:�7��U��D�-Z���y��įiZ�ӳ�45n�K@�+����S0N���:7�o8nܶ�NB2�֤a�ӈ�����`�a�uR��'-�di�Q��{Ǥ�B6����h'E@��ZUJq~T:��ăiZ�. �⸢��i��h/D�����Α+ŝw�$�q�P�M�C�Sݶ��/r-k�{hn�#�����S���%*��s���&�踘C��4~P^��C�8>�]�s��^F|O]�s.��͚�	.,�
-��+\�V9Y4�r6
������l�B��˓Kj,z^�4�Gr$�5�'ZF#�ΐMD`QS�����G��%]D:]h�<%�70[��OQ�Qݦ^�&���z��k�[�n?U�, �7d�wl�[�SC~W�m����̗�F��A�~�\�j!��	��ߊ��%�!A1Ė	U[��F=LL%�,�E@��!�T��@�׍J��>�������˜4\�-�g	!�jG� ��ƣi%d<�֊��v&�2U��-�|4�-8_���h���z��>H��+QfO:JU?��I������THL�^��&!��:T��-�U���� ŷ�?��>e���JAf(�/<3�p3ª�zg$���9XdzB�z���wY�o'=��%Wt��~㽎겾����z#����$��{�S��6�����z����
���9�5�.�Oߍy���(A�
��s����,����� ����i�|�Z�Mq��U�v¦y�D�6������s;&�%-�0ۘq ��i�t _ d�g�7�CA�O�Td
9���}\3��z?�ia|�$�����){lʅ{D]��.A�4��L��7.�5�1���w���e	�BATG
.Cn����!h��D������eWsջ��5"n
�H�&��-D��\"��Ժ��T��3s�p��*b}�v�v2�{�W�(4�/q�s+�'���6k� �����#���G(FY��&}$F��q�j�1w�fY���k�&��fLg9q3�~$�ms����;��+K��a�}�w�[�n�/ ��B �����k˯E�:;/��$�<y�:\���nx�]��BQ$�8v�13�һ�4K�V[�����b�[��#�o1I_9�%��r�{ЂI�T�D�z�H~`� ����&������#�J5�FN2{�OJ����#�]:�xy1w����s��`��@Ga�����/�'pE�`��ػ-�PU�3���l���Ȭ���$���Y"pP��շW��{���O�ޱ.b�f&1�/Z��Wg<�k�� ̈n�C��7V�r�E/;ʤ���.<�c��uk �~#���*2�q5��oǘ����#!��\`SP�Ȯ)�55(}r�l��&������ �,�y�y@,�����m�f��񸦒�V[ؙ��❏�u�= M=1�aeX�PK�pv��|/�����8�2z�fhl�������%*��D��ʉ���V�3FJ�9�+��l2�{�f��a|wCm$��}�a�� �@_?��gD׻�B(eӕ��?�6�)�Pʵ�h��\<#dK����\�v��:��U"+g�,�M������o���~�"�go�<�g?�2Prh�)]�Yk�}c!�2l��m\���
.�ޖ���cN@�G�xMԗ�w�|&�!�Rh�u��Qd�|ӎn`����{�b�*�r4F�2�$��nL�����P!�;v?P�Jt�Ĳ�֟���4J��1L��9&��M���h�2��iȁb ;������ �ᯯ.��I�e��c���T�y��v4���}��A��� �V̉������з��4��$xo�z�0��"��X7��w��}�(b���be&gb�cL��\��ڍ��aG�wx�*�qwd���	���n�^/.)C����-�a*��O$Rf�@�J��:��E�!AIí�Jd��+���.��;��+��ZL2�>�ʴh�f0[����+Z��B-��wڋc�*��'�c���#���+���\�kN"0�#��u~i�'�e<��C�C+J�#�Ù��6A��9�d��J+�ٺ����e��y���H��c�TЛ�9>r����D���jh"��@˦��p9Ϩ�3��]cq��;s^��k�J�B�#��]1���&iD7�6P�AY*��l�&]��#~H��g�6�Ƚ[x�`��	0��- 0JF������$������z�ٛ�cX���-�|��F~�u�,C��/�P�{n/b`uD������Do���	�g��!�_r��o���f�m^)�n�]��+����	sgH�����]OqIdҬ͘#-t�]�"�-��άܐ;|Y�:+�j�fn��9BG��,į�ĈO���{�*�D-�����k�����B�iѬ8(���R]|*3��i\�J��!^|�`ˉ�H"[�T��xIc�9�r�ש9�a��Q�2tw��auSi �.�W��7'�ɭՃ}qL}Ӎ��lc����qhU�#�r��;"�a�@suЍ�v��n �U��&�gұ��*j�F����BA���w����F�mVE3�ީ��Wz-��(�Yv��[yHV)��r6���#]W�gC\etFAѳ2��?�vj�)�H�Z���^�F鍌�Y.&~[k��b�P�������DЬ���#|}�O��ev�g`�d3�P?npv4m+�|��/+���L�7)�Y6�3��=��)誌��3a�u�c5R�d��m�5���.���`'H�4����T�z�Tn�Yk�4�6���J�� �}
�i����"�4NCZ��Ò�`���%�R��1(f���ul��u������Rp��.�!����rsΐ�)H�3~ȷ�W�I��^P�8<UR���R��c�	č��D���4pVj��D�2���-~�9�i�l[b.*�M���~��YH� ��h��$��І�FC��G�Z���wÜ���1�;�Ր�� "��t����B75{��*�H��<�sR�Əs�*�ГO�`&������=�>�P_�8�ڕ��X���V�Z򸾭�	n���կy 6l.ý=���i� bf_V}!�Glw��x�W7�c�4���ɫ�C��u�!�I'�6�
\��S�{�wC��C�~�9�d��wQ����pJ��8zc=�-��z���� ���\*j����?���|Ey���O�&	�/U@4�1�x&�A�8M��^�X�rw
;.!��˷�(�B'_��
"dY��T�j4�)��_{w�o���yzj�	��0��<�$��7Dy�h���I� �W�?���4^A�	�f¼u��5���f��"��-gZ��KpT-����+$��؁��l���-���:�Di>lji��B���H8����O�p�E_s����
4�}�>�`��0�x�����
�-|P���qOC��:���S=�A��_�fm��Tҋ^��Hf㩖,��n�=�&P԰:�C ��hM]kh�A��\����B�
��Dz�,� ��@=�ci/��!N�K�ʪ�z���ԯ�	>�T�!���N�_4j ���EkJ� :�~��C�>�8���Ͼi��'��VH}8����>c��Kt�i�K߶̿��ӕa���>�<fQsC7q+K�&j��O��t�ӹw}�����%A�~����1t�i϶W�f��_,��!0������n&��P"�qǣa��u���рV��|�(fd���&DZH�O{�pٚ�������!ۙ��{�@j���d��zW��s=c�Z���Zk��{�� ����d���4�7ɤ��{º�A�I�k��Q�y���f�v���O�_�d�ՈU'��jdg�cz�b������b��6kz"vĀalX�Yk��[%6�ˀv/fRa� gf���ߐ��������t�	C�4��,�^6�8K�@"�Lh����}@Ӳ�����*���t.�ω|�@��{fs5����WDF�;���X�߬,��6�������d3T��ھ�l6r3����=�L�͙�1��N�a�c'&&g�h'H�y��MI;�\Zk<�?���BJHKq��hۺ�s����]�sQ�b��iAw�?ݑ�����B�xq/�y�RyZ,+->v��?g� �]� I Wk{����:8$o�%�A��ulލ/�'dB�D��Q�'�\	��*~�+Z1��=3�dy9��l������VF����?g���3���W�ͳ{ݩ0�����u��@�,�A����a��V���0mo7 A�;ǹ�ݣ����Wݵ����O�Xn�;�D���֚��/��6��uo�"�U���m�%ʝ#� �Dpd�]�O��Qǥ��!�����c,j�|M8@4��3�0�+[k(�O�j	NT��z,��{|��a��7�J�2a����r��2I#&5���m�7cS���	D$G�3N _�����%c`6�e�ad�F�hxO���JU�@�cG'��x3j;
.��E .��BOhiJt'���o�(/��,D�>����2����E������ l�ܱcQ�^Rh:ԁH[nj�(�tΕ������egA�0T�s�@����4/0��h���4"\�7�=f���Im�#�w���cLw�V�A�#h$�7-�EC��3��Db����Y���n���
Z���i6v��^NJ�^/����WN�TG�]���&i�t���Su�W�5X����:�Z|�5ƻ%�Լ�Eu��y	 ��=oD�9�gzb�q�g����d;@�\�^��F��x
�-X�{m!"I�aێ���+��C�bs5�Kx����S��پ��4J���ߥ!��E~�;y6D�o�]^Թ�*$Z-�Z'��p��/�>KoU&�=����kp�^����L?	�
�z�"�R@Eo�À~���{��.uTUOf�4�,;�:TB߼�rK��>�����Y����#GV��Y��*��>=�G~'3_]*��pퟒ�N��2N�Q9M���N6�=�@"�OB<aŝ �G��ߞI�S �@�2��JRXO-�� ��K 
xӕG�� \tyd��v�&5k�Z��
�<�A/�f�ק�³�����F�T���X8O���W�6T�Α���8�w�@��_f��93OPSŉe���L�Ȁ���
Th��­��<�`��	pD��������ѳ1�9R|?��)�\�B�9�_�ݭM]�5���PP��Wػ�@W�U����)lz�苰� (�}�-8~sF�p�fk�BdLr����Q}�'|������j��*�+QZ����Vi�`�@<R�=q�~Å+c��~�"�GT�s�u��*�o&-h�y������z�V�f�"k`!��9�=>��Ôa�(�-ł�/:�J�֬ ld���z^�f��&xл��cN=��ƣ\2=�9#|V�pr�fc�@�	?����
 pM��Dz1a%#�,%��H�Ν7Ϝ�qt���ت<8�
�������(+��O6�>�9(x1-T�����P�����}C/>a��-3�.�%�*��NI��¢���9Ǣ�o��pd}u4��Y6қ�/�.�$xX�G�;O�̴�O� �{@�t?���z������C&��e�����?�]O���!F^��O7�x}�66�,@#����xw,s�������q���~��(,��ԭENE>�t?�jQ�O��eZ��3X(�Lu�mSޛ��.��!S�J�0�����}����܊\8r�.I�Z#��%��>�����u/:mb�:�����[� �ܵ]!e�E�Y��ȐM���R�d������Z!��d�/R$���,"��/��9�[$��	�=[?���Y�h�i�O���3�0�(;�c���A�7x}� ���n����='w2�y�5fk�J�z�fD�&��,���-�6���d(7a`S�^���*�s}�׻M�ؽ����s�q�7���c%�����C�Y�1����
��-�b���L8����2�3�Tͩ.-����A�����x�rQZ1� �9�R�1=Y��Ɂ��gI�@���x�F��sJ��A9K���ߖ�D�"<:i�Z���l��!P�ݢ��r��M|��&�uGe,���0�����WB�;SVV����x�z��l�]w���F���Ηp�A��_��\ujɬt&s�{�^!����A�ݔ��ǆ	�mT���3H�EN��?۠���5�Vn�K�Hu�2\����o�e@��/����]֍땍�O��*l<��Gr�e0<�'�\�����RO�� g��}>b@���@�aC��`���O�X��W�	��NO�������d�jByz;��K`��1�di�uh��5{�G鏁U-/Ld�6�w�CX���oƣU*}���B�G���Ǭ �&�'U�	���qf�>	���jJ��0����op4ޛ�H��O/;�MW	��&t�<J!�`���՚�����BL9<���0Q���]�|�vf��������wg�r�y6����^o��t76���,�@��,~�~�f��h���²C���l���S�Q�J�L0�.�O�Y����;�T��d�tӗ��c\�,���k�v2�^���,8о�E	<޺Jv��$e p��r���K&�ܬ�z1R�x���Ѽ@T�oni7�[r{j���m�T�QU٧)�;l�
HУ��j@KF9=^<,gz<�}�s�۳[�dMܺ}4UN��g. 
X�	,f�@�C����svB�!n�%�r����d�[�!ӘAsޟw���vp,���+���wU�Z��_��g.��s�0�%��!Ǹ�����f).*���f�i?��C�Jk ��g�ުI8�	�@�{��0�?	WV
�)�L���I�#�H�= ���)�p" Y����j�:e���*��	�0���7�fA���H���E��ɰ�C��B6u�!�	kF�����f@$��!N��(GY>tt�h:�2�@'.��=	��'�\u�<��1f�(N����$�1�)��%��I24�W���E�o��d˥���atÈ�g5Z.8qm��Ԋ~|7P�"��LF�	1���+�2전�GY�ƥ	w,&�Sڏ�E7א�E����ZU�;a ]������a4��8�h��c���r�-`n��ԓ�Q(�ˑ�"X�a 6ƛ\	d�S��=>o�:��F˾e=`��;g�"�?�'`�H+M�!�`��n��<�O���0�3�%�Å37q��:9�-�]�+it�*��E?C�6�T�֊���-�iB������SL����z��#2��3g�z�u��1�kz��zXL�J8V�Xo3���}M�f�/�	�O����8'�Dsx~�b���e+ԙ�?[�^�������r��ƘmKi@B	�R�:K3b����˜�g�6���|@��_^��Ut�\2���ix�՞p�'���[��:�4�X�3�.�Ǒ᭾["�[�^���H뾔 Ϛ��Z�re�/XR�掼�~�r�#������6Kq�#@�ӓ�Ķ���^&��&_�[U}�_ӗ��s�$��_|́9�w��|��m��i�r)?VRȵLe]ߣ���Z�ʒ�4�a�P �1s���K�:�	��^s?m1��ohB9�?���u�N	ݹbv���Ke+wI�U"H=�O]K��
�����~ $3J*yi��'�
����>��
7�)V��95��+��D�j0��tJ����Ǻ�Jum���3�ۨ�B&c�/�����l�ޥrb{d�<2!x��/v}�Bo١us_��k'*�+Ǒ����l~�����Ț����F{&f?X�е�x�t0b��U�̰8m
.ER'̈=^bC��dm$�T3@�����x���_�\[<�����������L�W�o-��$K�ǩoP<w,<���iۍTd���0Z�d�Yͷ�S��C��g��4Q�>�mx=b�|դ�t1s\�w��1R46�e���J�^��3^��UGcj��dC���'�\F�U���{��nJ�9�݌�z�����IU��9����@9O	?/�+�dܿ�u!�h)��fc��`;SW0>p���:싀|#_AW;ؓJoy-f"�$�G��m����d����-j�����}�sI�ܨrj�/�僩Xd��`Jc\
rN祟#�*���콕�<�N�ؿ��22��3��Z�|��ߴ��8B;?օ�,%X�;�I���hs.<���,�>�c3u��PԔJ<z��}�өb��K��2Z�W�{C�GBFe!A����9�nā�i��!{Czじ�2�CFU*=kO���U@q] ��|3,#Dbºx�{3�	��;I����5,��BFsZ��S���a�֡9����-Q^f����#���^�p�����g��z��!Zi���,����g��A�
}d�����(!�m�0°�[w����� z��´źC�=.��$
=VV�ӑ��wd]���a���\���l�����@�Dk��j�?��p2	EZ����_V�3���~E��������>����%��]��d[�������xmIS 6 ���/�lxSS?���qE�N�㛇C#����co���ެ�ه.3
*��iy�L�S1'�r0o��Mb�J����Ǚ�X��:���q�Q�	�� �N��i%�B��M�㔒MT�̹��s>?d5���_��3>H�&����R����5'V�K��P|С�U��+O�����l�8�F�ǉ-�7R5T�j�]�I ��B�!t{Ǌ3f��m�on�+�m�J�b��>e�R��ICM	2�@�{B��L~��_�vX|h�%2rN�
��+WQi��֥�ԝ�
t���|{���&�*B�f��%��4���8� ����Q'���-�p�c�4��O�;9��2��m֪�,*�7����o��� ^���b�@�&��7����&<�[彡�ap�i�ǉ4"�i^���o@��L��`֯*����K
8�߿��fQ��ġ"��<.F�N�Gk+�)iB߇��j�/�vp=)���4.)��V�P�x���IJ��ղ8"�*��l?���hjw�ΰ���U �%�wSd#ha :�ՠ����4.��v�:{�u�WH^:�\El�G5k�%��11@�R���[O��b5�/G�wP� �e$E����IJe�G�9��^nE�Np�`�������t�� +�h���p�{��Q&Kj���f�q����
S`�3)��)�{lP���!C�C�L�Jz o�!YmX�'�yS�];��^y�BO�e�:���=��a|5ZG���7_��/��^M����T���|�V%f�;QZ��K|��߰�����DG2;͌�{<�u�>^�hZ�
�(�Ā���Q?ΆZpv�^���g��,�X�R��&l��o6�9 ��l"��.K􇘔`�/X��G����~�j%��&����<�1��{ˬ#Ƅ8��M2��@ATx�J��J��iLSn�[63�����~D��H��p�ϣ>\�����߲3���������Dć�Y۠%ۧɼ�kv��k�p�3b��3��&���Joe���X���1(�L��,�;��j���9���� �#��vh�����%_��{�8�,R�7��ɟ�uh��;<a���o �CAqK!K@CX�_/AIp�,`3��*�F��W��e�ܪ���!��x���ۧ�-�y��
j]:Re��[S7�Ft��<��">��l�����|�B������/�W�Ղ1�"�`�2�Z^<�Y�75B�nE��,�H�U;��j �g�b�M�Ee�ù��jw)����w��6M|!2a6f*�֋�Ռ{|E1#'lQ�Ս5&~�{�L���>�������eU��/z��ž$sr��@��FC�;� 0j�L�N²V�,�~�"Rc�m����!(�49�˶4k�@�W3Q��#3�:�F��U"��
�5�Mp.K�{G=�,[+��W�W<5��E �{hHU.ҹK��d�����|�܉Ǉ�:.����%�p!l�4�����V�Q��ލ[�N_�+�oHrn���L�3�|~�d��q7�j~��a��e�Lq���,t�y�eEZ��)��p�R�pF�09{����#.����u[[`��N �W]B~^�D-����_��"^;����F)��X�����3W�ᔌ|��[�ƲDè�E��}�Ǹ��6f�8G��4|BQ*�[�j�.в�U���nś�#�Y�o^^�#��ME�)�aa���2ˀ���tZŃ�R+��f����񭌂��ʿ"���j�긥����,�e��&����,�	��|��5�u[*�})��a6�s c�G����%j\�-��S�a��&5��;�q����`�Ps�3w����(BѫP�p���&���I7����p�<M�A�;Z�\%���H��ݾ$��byC�y�'��x���)b~B(
�!�{��QP�.ԠPy��K56����Æ��V�����!�JB��-,Fqݶ�3џ��M���V���O��ݕ�6ŮrZi��p�<p+��/K�(U h��ՔMh�dc�E��V�s6u�E�	]R�`�I�:cƋ��#5�D��p����U��{��	:mJ��C�̊��ʳ��UBH�	6u>��T���s�筼���+���W�6��=m�����I��i^�,���*�"(� �����:)K�-�fɏr�(P�\M��Z���e@&#q$�fn�1�!���W�5'�+�����K6�*��`:!��*�ىt� ��S�uP&�ｗ�_v� P�I�#����<|	%��1��A�J׍y�9�l����-�&����q�SE����7 M��Z����1Z��K�����j&:�Y՘�4�Ù2'�on�L7�.7zv(�bܪ^P&��w����)
�>�%Va�� ߼����;���^�"0�Z���X=Y��I�����y�R�#�,05ꀹ�p�p�JO��1 �\u���WI�,�U�Df3ڴA+��P�).hz̉��̘�F;�ߎ��h������W�#�jJ}�2knd �K	��u�%���Ss�Qn�UI��V�C��w�|��׽����
�7+����?�t:�3�)���V���� �=�Ks�BL=C|h�~�s���9z��+�e�/P�$�+Jj(2�e���z��oC��j�*2ߞr�h�I~a�u�A1��Dt�6�B�8�&���s�(�2�MW��C�2�l�(�i./���=>�X2��w�_�6h\_-CN3\�ŜX��hϺ��<Øނ�m,�������� �(�
D�W/����%֟0d��߭A0�T �#Ex|��Ϣ#o!cA�L����rEY�pj��AU�x�7�%��K�����3�k���m�&�m����;ګ�+Y%�Ɔ���?�����# ����<�~OY���7Q^"��]=�!J��@B,EOYr�B_����sZ� P(#��
��$�{����庶�}��ʾ�/8�u��qV�������6Յ��^��������_��q��>����c/��U@�W=)p�4R:h��{���Xq�g�7���|�Ӫ���B�E;�A�\8���xQ��H�g-�h�L��'�U"�vJ(U/L���h�`��$���7������~��>	�Uf��)u\I$��!zk�a�G����V�d�<а�\�ia��1���y�njV�>+��*���+�a��m�l�/F �vah�=�0M��gK���~��v�j����A�v�-D�J.?�o��.uD�C-��B�'�z�˾�i�4�/��a�ǐ{1̜�@���T�U��%xKx�t���T��+d�uW��H 9WQ,�K�fu�K��f.���տU<j�_�A�ت����{�/�u��|F�w0���.�tv�fs���}����;�"0� ���ka_��~Y �����S���`����M- �lR��u1KD��򤤁��S5�%E:ߺK9�,S�����8�?�"�"Gл���aQ.h��0�M��s����s�ޤ��dB�<�����y��lb�kR�k�]���	lL�2�6�Bp���b���=s�K��}�x��w�1��{Hf�
����x=�����Z1��]6$�&�Z��C�y�]Y�H׼xo�=�����8�Q�=��y�.Tˬq�f=��T���mn�F����IF��j`%OPF��K�E�#Y[�g`�I�j��Ҙ|JZ�4֨=�I��8���� m���Zߥ� �
�x��L�R�Y��_�4�f@畵�|3龴r�
���C�oHQbKw�u.$����;Mw�NV6˜C�����hbH� _£n��i�,�*Y�!FIb4�\C���C������F�.�w;)
F�����*ߐ|o�*q��Fi��M<�Q�0�����/�Md���D���Zw�z<�ۜx�����
���_�lf��W����y��v/��|Ͼ�����rc�X���.�O*A�������CI���j��Xr����H���I����t�K��?B)�^~^����֚�T^8X�󡅶e(���<��C�� ���kHTa��jQ˩����`��F ��2A�O������[i� �9�2�/Sr�u�^3y���T�γ��̛c0e@�"z���ٕ L�殅��h�`�-�B���=��}�or��e�� +��&GST�oyl��x�nҚ~���&Aپ F��dl��V�����VUO	4��,y�U��Ϟr��Y�ñ�[.�WQ0D����Q��H�O��
���g�\<H��)%��� �h�f���_滊��w�]���n:U�ADtx�p	�����{#��P�L�xi�l�"'S��)�JQ_���]r����Q�F���K�]��v�	@	x���x�H ��n �|�|�n�KfT�Y%`�Z}@�v&	�42�ɨ���4�S>�`�姄�r��h�N��U� �Ea��	�M��I�̜W��̊���NʶL{~�8K�ف��Ͷ�+Qt$@�땾z�g�EP����O駰����$�u��6*OH[b�+�g}�&!b���N�i-�S`_��(���|)��X�7`,(�~7QUI�v�\q���T�4V�j�7`��p%��gֹ3lSբ?	w?�Z�|4Ք��!��b�^�^Q���]dA��$�,���=DB��@��3����*z\�-�B�p/�bU�c���Hl.&@x��jQZ�;�0O_f��ꖥGʰ-�6�h1\P~
H�k 5��a���و�oIa��{PG��(�jD-<���1�5@�؃���y�w����MCԀT�`�`O�	�X/8�Os�����f�!��^>��;�h_
�Pp�z�Im���L��H)S��8�m��`��d�A�wˣ@8z�r�0�q?�-&�D����"3s�?7�L��睈�d�ĵs �x-��2[��׆t��.��"QcI�ESzSצG�Qi�.��v|��ۆ?Λ�Ǆ�G�	�,o� /�|��}6���Ç'"�R����+�҇��~���Y�G!�G�u�����vCs
P�)���A�a��$�1,� ������FZB����$��a�7��Z��+Q���@pB���	A�T����;a��Y�)>�Z�8�)~Bx�P1��-�n�S1)NG����Mt�pL�y�h<�꫋����QN��m���v9�E���>��G8�K�h�G�!y���v=�ϯ�v��AJ�	���d�w�w�4��
����V=<*1X88�r�<��@��Oq K��h�/h$��ԝ266J?>hq{JMV�m.7��l�F���������Լ/mf#J 8��8
V�=��	����l��.3jg?E�Β(�z�-�&��>�q�iv�wGG�ﱏ�B��}��{�~�_3\�W���h��\
t�.���]~��_�յI=�eM$Q.�Z�q+������t�b���=�ȋ�f������(� p�K4��+���7_.�A|5WLf�A���}ѱ\'���9`Q�t��SꂵJd��nv����ol�����/�c=�n���?5&Љ�N�x>���ot�ߙ��>P�ȷ�D�J4�޿8�%��Έ�Z�J.����P��D���5a8͊)@q"����1
A���C���w�Ȭ��C����6/c�-�]�`wT�S	{���y�X���T�A���\u��;r�&I����|�^{-�D7�9qH�|?��:JWD,�|g{q�35L~���CI��+"�[cK��y�'����pqR2P��(}�����y�|Nw7�@SP���v��\�Z�?؀���l|r�.��^�엵�҆ی۝)?���=x���~�de�JL���":A����瘚;A�H��Z�2��g(�0j�/ -�\o�c�s�P�G�O�`iX����Q�\��_���rp����5�#�f���C�&OM-��Rs5k�Hy
��%���z��l�kY2��ۘ$��@���/5k=�O�ϙ���-	>9Q���S�('([Rv�*�Z���ȯV���f���������q�s���w$�y.���aX�8e*s��Y����[�6A���I���`��O@,�̦��h�C/��g�|�X���l]��\�bL;"�}�^�U �}=���
�}�+h׷66�mFE"�/�d&5��z�c��g-���SS���e	���:39�<-n��zp�����9ڨ��K�Z=89�/�wz������Z�b�����t����a�0��q��p7�?�����L���lޢ�B�������w�Wm�Jm�y�>*�����i���M�c%E�y{��k⪌�}W ܮ@�����/�}�u�f��ȉnߔr��ڹ	�עM���'�ʳa��8A�ɬ�H��.�@Y�C�;�(��rk�pc浇����a~=:-�_n�VB�n�-^������x��ЫV�yJ/w��Y&;B�ϐ�a�}}�b��/y~T��G�SC�hӌ ��xB�l�Iɫ� ��T�	��9�ʂ9�'�۽f�'_�o����몬F�W��c&���r��2Xݕ�|j*q�ڠ*����u��E��Q�InJ��8[��A,�"�UZ�~L's��a�[r���V�Q1���fE���X�⁋�uu�d�2z�@�w�޾���?j��T��}m�'�#��N`)i�Z��qw�78^[=9���yTp�L~�F{�K��T�O;��ʝ2��b�9���p��(�5*wm����z�Av`���B��m���Ə�I�ϡ6���j�- ��|C���o>����/q�Mk0�Gd;����Ҳ,M��Y���3VI��M�hBJ�E
ĕ�8����^d49߆��8a|�K��/*�w�ñ�ÉTF+DxBM4��}�uPy����.%no�_���ּƝ��e�}�0��.���wձs���U�ex���$D�y�CH#d#ȲD��;c �^�x� 4�Gq0�1��15����A�\�! �~��?:�X[�+n�y���^M�'�V9���[�=3�\��z���ۨX��[�s��v����8VH@ll�Q�7-J�U��� [zt����MN9��h>��sf�+���x�柎�'l��$��3�Rp;�_${��)4T�L��I�%�Bְ�z�*@l�Bh��C�Z(x�1pR>p,u,\��趦bD�_Ķjע�0��*��X�|Xx�>g�%�h(WT%�e�Vu]c�{q��wL�������Ro��1ǝ���|�h�}T·Q��aՔ� �9��nq�4��֖I���
+yr�s0��4�;��.1������ʤ�r����c$ �#U2��l	����	�VN��͇��X�O�yLvkb�Z� X���8��b�ƒa��.��GQT�X�Z�Z�vyE�m�X.5:Y��4�KEIG��D��G���A�u�z-��h�/XPz#�P=M
w�Q�a�?S���i��5Q���G�jJa�Χc�m�NM��ݭ�ƌs���jg����5n��^H�<�&]F�1����)Kr���%�eU�%NI��dn��)�ktt�v��h�@��(3���cYh��qO6n{O]Kv1Dlh0��J�&�!�[�N���<tb�=����'hP����Sd|�����1~9���S�#O�y_����j�+x?��9@,S�(��`��&ӓ߼|z��� )�V���Z}��v�̩1m�u�r����I���>�2c�������|�	�Byb�稳�#��,��Q����?�k���Ʌ�A��hC����c�n��D�"�̼<+lÉ�鰆�G�"�=5`~��t)�/�ɻH���61�N�-mi��z�)K�mQ��-n�ӶYDf�KEt�_njPB>��
V�����L�r���`�"�e�[�|k�����ADo��-��̫vt<�\�[����nCh	v��@�Kλ!vn�<B>(C���x#".��>�����xs�I޶ʥ�-~n�A&��^D+TÇR�0d�7��,pO_�o��yZXW
c�s�L3#��P��H�Zt�SK���+9�X�2���Ƃ��jd�{������_v�*��ȸ���Y��hh:���s
b�T�_�o��X�Ʈ8$i�Sw�q���C��K�Dݞ��]ܯby���Qw�I:�!���x�H�-����W�`�������h�&���g�;N����g mHz$�8zM� ����9�><�.����X�V�z�d5����*�rB`�1�rp:K�<wOhQ��ծ%yME�&	~��϶���;8;�p�OF�qzF)��p'��p�y�r½���*��	J��*q�4�/����/�g��C<$J�U��-���;G��O`������V�5$��dn0ѥģ�� ?C�m�D�	3�ِ Q|���ߪp�0[gE1�Q��$�v�8�/��(��RZb`Cg:"�N��휁�+�Ng�r���Ӭ+�X0�t�-�N�|���?�
C�� �L�^:n?�+nڿ���>ƦW	管���u�вX�|��tN�s����J�BC����-�����]��n�6W�΂����i`�������F{]�x@�7�