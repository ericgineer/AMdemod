��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�Jɰ��^Ț���7����or��c{��E4��S|7�l���f8��r!�ߥf��=0<�O?��F�*z�������!��v�����"}*4"�8����:x�nM�,����5��p��TK�����ހ������̻���ߑ�*��Q0V��q�e�gڇ�=p��~��9�K�Ie�����/��ȏ�})�ʈ.
��i��}�R>o6�3��D�!��oܝ��G��'�I��w�N5&����XN�Ycdf�AB�2�ϑ���a����MҮ/P)�S<�>���T��$G��������<G��V�������d�� �0�#Jb����O����P�)�̚O�r|ɪ��5R����w�s�h�Yl7B�|,`|χn�T�E��/������3�m�l/�����/I���Mئ'K�̽tVu_j({)s���I���,�f�&b��|�k!�*ɲa�P��RZ��D.y�")�G��W3&B:qP�_8t.8@>%���:�UU�&�HCaY�j�m�Iݞ�]	)��Q|�z�J2�m��*܆\�<c�� �� ��]�ECw�C0%nM� �G��Z�RaێM�$Ṛ�ig���^�S3l�d�������ح�����i>�n���������y�;�l�ld'Jڻ���B�5�U��F�*�w�.9TM0.��Jr�P�>C�RY$�sz^Sl"PB��-9/ ��mT�È�`�c��Z�]�
X���܉�y9��y)V��L\�̌D�o���bEt
��P�(�&��t�B���L���Ξ��$�Vቘ�p6Y��ƶ�}N@(�ve��M@�CQG�� t��	a���Hd;�JJ�D��l�H���bx*�ML ��)R�&�۔v@0y�Jg��w	yeQ�4�ON�o�Y��ʐ_����MW�g��q6y�RP>��O����nN~Z#w��!%V|X��y��Df|(���N1WN췹ٔ�[��	����Ip)� ��������:���܅����b�I�IN��w
�"�������5K3Y�e�������f$�Ci��2�R�35��/��Ӌ���P�mr�d�$0����)�2a/�tP~|E�}���� [w�ӕy��;g�!Z^�"���޶k��
3��ߡ6Z\�T)ǫq���I(�v��5�rTWd�U`C��XF��3ԐTi���?{��*t�C�^����@ԙ�'c쮜�}������v��됊�O�r<�Y�i��h�����-���\���T�b!i�c��5��֙
1J�"��e�� �~�L7
�id��J�Z��t���]^e#+̧�[䱡S�)����k���X�Zmd���1�f!7�������[NE�Lbe�"��[9Y%�@n�[Oѩ�����\~!-5ȷ�������}��FW�� ���d��'B�