��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�4��~�4���֮�+��o�6 k��ˤ!�4+B��rx%��s���`��g'�W���U4���_�U�:��@9k�|�?r7_�����^�m�4��6��C����Zk���z��)���u��l�ͣ#:��"�ۛHB6S�=���8��)�PkX�cJ�}O�C;��0(�* b�u8�cH� ��,uVb����>}w�O*�n%L-0�t�i\�:����>nm
�Ȁ1�XXY��Rd_Z�hG�s�� ٽ	��(o�G�>l��2��4Z<�2(ig� �We�{�gB^��G5�ۧ��X��_����F��I[q�N����������N	��3��w<��/�/p_�1��E�w��b�����F�W�<l�#�iڝ�pt-�����׫�!yT�-~��T?W�� =��{I�Sm��˦L���4���.�e/1�v�9+�h�n��h$s�۝�8Z�k�ş=E��?�&�TZ��l"f��8�l�m��þ���.��S������JK�?D���YZ���Yc�Qb�-�X����#L�%B�3�r+�,�6��V�*�cե�E�貾�M���Ӕ�Y Ϙ��"�r�l{�n� �ma�!R�N��y`0�k���YC: �z�6��tćIz� �opm_���Ib����ʭ�j/c8W̖�$ph"��̐�c��L�\�H�2�Ob�ؒQ�p�oՍ��v��R����l���9j�i���k�U����J|q?f�������t�^��6�R- *��c��]�k�Y]7�tX�E���Y�q�u�Wp��F������0�[����}@���H��e<�]���;�=�Kq[/�/y#!�V�62�/���qh�R�۬k8�`$ �ޝ��M~ɰx�АRъK1���Dw��d�c�n�D�.X�ח�� W�Yv�h���#��5)z�2���dOǚ:Ư���-�H��P-�ߝl���R���f�I=�׾�+d�� �#N���a��%����-�_ѱnC�]�i��+�a� [�A��`��q{`c~�LT3(��PX�oU��H����M���V�r�A@�m>���F�؞(TI�n�^	[�[������@x�DI}��y��"\�,>Dv�=��0@č�FJ��[�P��MM`�ܶ:�.B|Zφ erе��Pj>�+���u�P�"�8EB(�f�ʖ̍;u��:Qļ?�5^Ƚ�,Lʟ]�F�G"���a�aIDJ�_(�[m}��`3&��X�K�-�u���ie��� �B�6w�±����NF��}m����Qf�2�UǷ��{��#��S��j��`5cJ�:"�LV5���{B"�g�)h�'m�+�(���l=K����}����e�����n�/U�l�% <�����c过�;qI�D��u��C�>2����c;���I��z���	� �M�'�<��� 3���D/���h^1���2 3��ґ��#>��S�Əf4���Y�� ۵�����
a;�>N�Hd�>�A�N�Y��I2X7ד�'�n��1\3�r�G��[L�d����m�`��r��?1L�.8���7� Q�F�mz4�g����V�&��4��]�T*��P�t闊��Hg}�i�Өh�B���%��P<�)��8C:̽7��k��;���?o�)+������0X��үWM4���.�hu~	��Pc��h�;��Q�B��Ycf�Ѣ��_�
�0!*���ۊ��t���"ֈ��Jɰ�ι����,Ͽ�I��2,�1�����c���d�6���Y��
��� E܁78ƒX�X�p��ͤ��O�WDpzK5��r�{. b�D�(r�v���l:6���Ċ	4�"���ХsR.�Tφ9]&�5倎!0��"�Vu�W�CxR��R�M���9�܄�`�����Ͼ!���X��z�<-���Ҧ��
6Ec�bt2�����T�|�(�1ߦ��6��3�}�z��|�ŚG��l�MJkF�a�+�5辥�j��ਯ6F�m��O<��V�B'mNC��dΟI��5�GG����,؁��TY6��C��o��Iv�ɷ��1Ā�j�F3�w��R��������ֺ\��,J KkB�}Ҋ�z�<*��b�ў��Q�5Aa_�cSϪf�n�6�@R��/��s�U�Vc��P�2NLi�f����)e��f{ q���m�����Rƚ�j��	9k��
������!�+qu���(�j����B����`cj>�ҝYDGH�̜�NZ��.g[�Y�g��:&�6H�v� m�msrY�����Bu���~H�b���6PF(l%am��H���N���$>��DXT��O= w������2���/���T{�>��^~
5�W��W�O�#N%9��E����w�v%d|?+�/��i����)8�_��ס�;z�MN�qG����:�O56{��0Ѵ���(��!~�8�3|��p`o�3[�V:#�Լ.2��Oݬ�Ӳ�V����PS,���uooR�/�T��U1�S֘�~���m�J���&�^�G��IϺ�J}Yy��*Գ�	��:�ON$p��wS��D��_S+$˱�e�aJH�o-H���f�}����*P��6��Qs�A�����/��(������.ܭ�aǰy�Ϭ��Ap7v��n��2�K�!I~���Q��'�5���⁑�g�߮�w�]�^<;02&�Wi��q�%�)�0G��/?��avAfJ#����ӵ:t�a�����e敎�!9uc�6C�&�5�Y���ek��I������+�b|)����*N�l��+��� ���ch��[����NE��1)���C��?