��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�O�5t�"��� ĸN�V�)Xq���!oA�㝣�V!��(r����6��DԓB�ee[�4���j#r٧a��������9��նwo6���6�"��ݿw�{,c�x���	��
`wgc���2�`t���o�(6Q�����w<�t��B�8�Q����/�=x����Y����q��Z���̒&��0Lx@��>OW��n����=r.����Oɳ #Y�r��˅s�jv�Un8�����^��� �5w�߈ Dä*f��4Z����YC�����'�z�3rCՌ���m_��'� D�^\27��l\1�H�v�����
|���r��?��yU�;>�*���}�
�GR}�(�h��q]O܎�)�@B�k�����<`�?�W풅��rW��l���=��P�û�$Al�����Xvޏ�ͭ-C��L���'R~��Z�bNUk���	&P�$�14FR�;���e�y0�Z5=�2N7)D?���b��M}�O�N�v1E"�C�M����Y�А�3KY��/?3T�{����9^������(l��~Cn��GƧ��d�g�T��9d~8|��IF�!qK�gk���kP�nѽ`��_�-b$	T���+g���C��M�r0D�I�t4aH�'����Lи/r���hQ�n��1���s&Y}E�G:s�O����9m�gj�j,z�}o�������R9�0 ?8Z��فdh=�}�	ǈ�w�	��]V��`�P�?�b:XNǔ�E�1���/b��nv�^�j2\����oiX����k�B"RU�5@i�׏'US���[pKvu2���2�z���Ǚ��R\r\�F��W< �@� L)���Wok�Z��~VA@�����MK�zz�c��>R��5��*��6����_μ�Պ�8��<ǜ��m7�f�pt�N�Kݝ�Ŏ�ȁA1~���Ζ׺g A�r��ɆHR�$I����EMt�)�Zq�׳��~͡k^h�Z�#䄞�
J��%��Aw�2'J]n�ʕ����aPTh~#Q�GOB7~}��|+B�?�Y*�k��w/Y�(��l��ۉ�e|!�bJC��HF�A���v�bO՟��F��~���C F�-e�� 
��G�\��&Y�DX������b��/g��@@��b��XYP��L�,?2c;�+D�l"yC��P����fz��9Y�8��I_�-�$�ANfy�?k��tn�l� "�a��M?�`}��۷1Dڛ�}go-P�+�Y���T��|��%����ĸ��Y�9'Z}6�55�`�2�і8�@\z:INv畡~�ޥ�u�㬔3B���B��Κ�={��
�s�?y%�w�U0@��'�b�}����4Bz?������L>�7c`d��S�j�S�kpH���;�D�<g������W�R'`������|�.�vit]G�H��M����o�o%z� �"p(t华rGSG��L�����_��ލOn^�Žy[��7�в�'' ��ʘ�=n-_l�y�rBK�&����>���q{	�'e���
C��ӕ�2e�!�{@�\f��Y5F�Q=���7q��c�� �&@e�8��6f�Y*"#X��0�~7�PJ��u�l��%)%��ʿ峊�4Q����]r$L^���`%X��I'�m�̥%(X��f�����I?�a_�z ����>�����L�UM�3&�O\�zy��%H�qz~��},�#ڃGw쐄���`� o���[�p��8Sa.ԅ&4�#�ª�S;*s�.1ŕ�X���404���9�Q:�����E�%�Po���v�� V[V ~�����$zi��O�A?���ٳ�7@漯Ql�0��Q�7�*gӺEe�q ��:�^�h1X�h���
���4�f��O��ه�+pQ��k�7�w�r{i��� �%�t_�S��7[o2�[ʲ�^�^��ƍR�����Ј-�<�2��F�p4�-�Ԃ�>2"Z���UTz��'��2��5���� ��}�J�1t�GXF6�
��e�y�余 ;_!7
����R��te�F~�:3���[��#Vp��Ψ���.M1�h��7�5������P�i��[���@u�*�
~���	�~Du�V���8,��,h��{�}m�YB�n=��rQ�%���5�jՀ��Q	�X��L
�R���*ڽ�n/
Q�T�"�X�d�M�Y�LW���$���<�y�[j{��,ʒj�A���ӂ�e!6����prox���H�T�%��F|�Fg˙`�&L��q��2���F�r�\٥�f1q\s��y�we!�L/��>}�8n����[QMQ�� ���n�WĲ���^��o�"UL��M�={��G�\��t!&�I�j��>s�*D�F�e�w�������Q���q;vڰ�]�UB\�p^~t�/�H�5��i�͔oAbj\�1 ��8X����v�K�Y��
	Q�L��Z;(�w�\mV!|�n" �IHm
�G��@�T�&A������R�\��x)������� EC�:Z�R[��_HkF� �'a�F�Ʌ�ԏ����n��4t�� �t[�?K����1y�2��M����$��#��(�oҡvZ�E=��:o�R3�8q8*��y�1y��3	��&���ĉ;�[lr��\�-�0��aQ,�� zc@뿦��߼��o;�����cWA?J/���0�3�/�P����Jiu��oF�v��Ψq���]�b�{�߾ߨY������պB�
t�����a<�)W�c�O���9���8����5�ϴ���ԧ:u�j�3�x�-9���e S�	*���搌��T
����0ޑW�F��D��5Q�wv=��M������3{����*��]�W�F�w=�/r�� _l 2���C~?�Y�!cq�a�Ěג�`��$c�8���~M��A���%�2��y��!a���}��+�p��c#�� ҥ��8�I�$s�=l5�5���Hۘk|���t�����$Z�?���;fI��S����V�?�S��1�H+�� \6XR�f�T���B㚌
��O��~F�ԣ5���%@i�I��PL���D����9��P�lN���C����k*ы����ӱMOJ�[(*\I�.��ֈ㫌c�ky}]���>�'��Fb%�̤���*�l�KI���K�\�éi^���^�?�@U?��)㨼p��YOr	�U�i�o)G���-@�E"O�k��<��1g���^0l��y�PH6�p�/��x�Ԁj�$���F�e�ɢ?׶�B�� �-��P�0��mn}�]��\%�U�\ǖJގbA���9ӆ�s��PW5�4�J�w�T�����w�՞�p��͢�&�����/,}�'h)��8��������.w0�/��i�l��c:�x��y�]�Ҟ���d�3�Ǿ���`�UB���7m�
���Q����A?k��!�
7o��ᄢT�!��]W�Zx��WYH��o{�^ҷzq\s�+���i��ip��D6�\�-a�<uXV@���tn���-QH�Rd
�)>�G�nGu�z�n�dYv��c?��$}�qTt��s�S��?<�n�.��DM��� �T{��F�,��X��C�l
9�@����p���o������C>���I�G�l��O1��p���dY�J��s�w2�r'.'t�����G9�[�'
�����+>2�ήP�\ (�"75b`,-5z�1�b�����%>0<wd�ƅ׋x��q�^��̧���C�~�~�z�u)t=�<]1��$'�-QT��K�Oå־�D���QK��/6��E�Cdi5�(��@�_�["��9�����$��o��
��0�iy�#S�}R#:Sn�A7��2�o�$�H��I٥������D��|�>5t`����O3,0m�����Q�t ɥv �B��>���>;�U�O�^ם��v�#/�{���l֌'�3*�+ޘs�m�S@5=�6�A S[�[�+څE�T���8Z	�=��a6��+�0!n"�r&�-v��M���1w-���%pݘ��ЫzK	.��y�*���Ŵ7��-��\��2L �~��UU&�I�p��'.٦�c�bs�j���.c����̑떲,P����&Օ�Hft����˔4>l�Z�r��F wg��I;�����=�.ʻr!'{ف�:�����~6ךAC2�K�z��XGZ�ʞis������f{g-<y,:%�(�5�{��.���Vh�#J/ ��J��ɽYk�s��O����I)�9��0��B�P<^���^�*��U��ŭ�����Z��d�>�0d��
����D�;�鐲�U���������ݷ-9�r�k�$)`��KZ��K��&���� ����W&���B�� i�Jב�&�/M�8�g������aE���hG�_�^����*"�D��ڞ$�E��^�F�k���Ӗ�L��=���� �w��5�����wbm~��Τ�'���<��b���K,�g}gU\��F��w�|	��V���i��.��A��t ��蘨;�i���}sM�x��92L��t�?>��֚�J3RZ�4+�ć�t+A��Ft����m��U�x���8�E˓Ŕ���c����pRίL��fv�������!���Us��Z���?ϥ�������ˠ;u����L�*�d�1�҈Y-�1���xWkŅ&$j����1�Q���0�)��5��Z�["I�	(�)
V+\�Dϑ�1�1^1��7l��R�ݔ ������'&~����O+7�y�Cl���~���j��0ŕ@C �^}�\bN� ���,����S�X�.D����<P�#�Bb�/\�מy<�Az�#��X5�������y]��|<��>Df���Z4a�9־��)�	��˶�#}H�>b�@�󣖓\�f��T��C�̋C�������(S��obu_:NQ�;A��
�cY�"to(_��7�V�kJ��D�T9���.[F^��'}��J��S����6��|�_�'�W��rf0�儉x(�j�Z2:��~�,��͸K6�`#t\��{�*k�KƼ�`F���U���G���������S
��:nO+E'I�Ǹ����R�u{S�4̻?��������n7��`��ҙ���h����F�n�a(�W�m�b�3�;qңm5��ej!S�i�Z�w3ث���B̻���`�o�bŇ�|<Q���$��ɬd�
M�]%��ɦl�/K��8�AaO�W�Y��^�F��7��hC�{E��)q*��c�H)G)hL,�5���Eð����f"o��,��,�qD��me$t��;��7Ć��u�߮���.�Ck���d�o����+4�c����|�:��;�	�͕'XyqyWM�љ�����ˉ��(x�+��,l���N+�&Ñɋ<��#���%�ظT�K��8���q�N(�n�F��k�i����1������"�vevʦ��JU]��e�̗�紪�a�4q��I�y���B����ɺ}k�"EB�;�*�q٪hܮ�<f���v�bfE�5�׮��R4����������5�S�m�E�z�k}'O�k���=ؘ��Z�����|�=C�1���9�H��K��k����6���;����U�L���}5"���d���`m���N��G�-���f���SA[��l}�ǧ'QKy�E��9���7�\B���w�7��c=6��S+9?�������oZY#9wv������W�y�L�c�,��c���k�mo!)�|n������e/�6���J^oc|������zо�
���[h��J��B�w�8w��E0#/�6�|���&���!���N	��"H�|Cw��+܈wѥ|�~b����)�~�X?����#.��F:��N�� ��Y��f���;�ֳ���uU�L�MwG�x����R�m�-H�Ud�w���N����}�NAc(�_sF �X�i����C!c�ĥ OUr���Լ�sWk�65�/���,���u�P��X�!�.�iw��v)��6���i5:S2 H�]�G�6�{���:��q'ȮyV���Oy�]��H�c��<��n�Z�{��d�e����,��,!�cw�iP�~�&�b4Lq���c ��1�&��.f�}���$�X矶�5`}}Bw��;6T�^�ݓ*U8�n� �/��
�6<h#�_��s�1]!�G��֭j�u#Nn锈�Je����^8�?�ަ��mn]�Aa�H��=4��J��qLo�ή�#��]5��d>j�dQt��:=6�2"��+�P�q���w sk *�Z��%���X�:l��n���b�`��Ƌ�
UsҎ@�R5S���b-A�l3���'ϣ�2 �Ţg��h�#W��l$��+� �sb�G�8�4�`�T�U>"U�!��;�m�8�]F8�ۺzغ���/1�nPX�qBWV�����ܫ�jX��va�B���PZ=c�0|Ytv�ץ����1�q+�Q�{x���&�$�}���T��.�����Vƥ��R7���x��=eJ���D}�|�z��Cw�u>�&D����kWn���u�'�a�X��3|�2S0���Aap�"�Q�K��O��x��Z��Ec^���`=x�>�NgT���x��5s��8�>�L�(����^*n� 䑟U�2�S����G�(����=I�k P	�|��{@��&#<B�F�/��A��o���CU� ��5}�#E�.8w�a�j��aM4C���gT+���@�Ct��GΖ@J�����Ѡ�E9�o�d�a�L�^���gR��g���Y� U�~f[��9�����j��&B�ǋ�b��~�\�	Eq�%�F�m�T2�=�2�T����}#��$,����M�@��+õC�:�<Ն��y_t�6�I>]���}-R��S[���ш\cH��'�)P(E�L�>D	��=C���j3�6�&X���	�~5Q�֥�e0��w���n�f��1i�8�ÉhRy\KF`�z����8��~��|W8\���Ţ������jv��N����ߒ�]�>g�wOձ����|����F�jz ��_Q�79Yқd��EQF!�Eٖ���po�8/$��T��4sHp1�'"�`�8����G�������~��S�`�yt��h8Xr��N���ϹD':��T������S�7=m.��s(��DZ`�]c��,Aϲ��������HC�� ���~!��ْ;����g���|٬��X-�N"Wǔ���xK3��[���s#Æ'��3�L�`"W��g�LәRq\ n/Oqi�>������ϗf���yg����n�����Y��ZӐy��_� ��h��{=.˰Q��xEYQdol��,9S�!��� [��'W`�v�m(5�?���&N]gO�7����&*�h�:( 0�(���;[��y�"��6���Q�`�%��X�G����G�wl��C��d��)�g�Wݸ����$=ǒhx��E�����n_�/�����ОO&���"��z�5>i^���K��wG�"�$��yt��� ��ϔ� �2J�3�Ci�JW�L�6G�qȩ���@�QZ��I��n:9t�a�^-F/+-��r��VYg�S��o/��Li&�X�p_��\R�n�A(��ja]0�E�	�nME�!���p�Z�|��<����YQ_�<S\NS��k���	���?N{wl�:��@M�ꅻ̧L��2��A�P�����u;ؾhU�zIL R+���wc:�~Aq7����'�(y{oeSڶ�l�R���mQE�-��8G1{E�}(���1��O�g��ȏ�����3���B����ㆡ ��3�8p����N�r���9��N8&� �+([LU���_��}�o��q���Le'��˝̈j`OSvf�m�d'Xkb*hUzt>�U�Z�$&^��bTi�Dɷ�-h�(�˽1�Ǧ[|gM>�Dr��O���~R�����J�M�k�� �ƢB���c�?�L��ר�G?�au��I�[���tR7@��\�T�pkj`�1	5~1?Bt<��6�����/�t^K-;h:k�"�n�����M~��5��ĠnB�̊N����T�*��pߕ��GXs77�L���
�5�.����@�zl}�Y�"�������~�C�DX�v>{�ƥ8�� ���+�� _����sys�b ��n%����;��*���yV���k��9�'U��m��[c<wX���t��U�hj�&�����E�z#a�͚��j^�q1�@�ު�U�v��Lۣ�4���
��z?�p"x:�	@�G��q`yZq£��l4F������j勢PV��F�K�3`C&�il��O(��Ud��)@g�͂�Cm^���'\�)�Z�\.TTpm�O�S}�J��B��Ύ�V�b�� �J�������yy�ۉ�T�����*�U?hG��:���&l��.��g����,M�K+��0��V�!����g�ݟ��'�]���ʽ��x�?����nV�L������eR�w��KEy�b)�^r�֨TR�)nU �u|�G����Q+��z�(�ݎ�B��1#P����0X\�a��6Z;����|�g���Ӊ�IM٤^��A���<�)?�&�7��")�ϫ��8u-��%  �p/B����X:'
��A�|Bgz,P��wt��:��	���;)ױ\j�;�W1@����q0\��l�ҟ�(T�H=�l�ԭ�~8\�$�J퉉֌ǕI��	Όz>��t�0��&fA-|��)�؆r@3�t��v�ѩ\t{r��g��b�N�c$��yL��}�0��f�7fH�-�b��� �k%�;�J���Ǹ�&c貜.w,i�����W�$>7����M�	�s���W�QO�<�}� �������j?.�R���+���I!�g��M�(�L��e����)|Z@���9wD/��H�L��}���-�YEyۮ��:��C�m>�C2��V�ćEd��C��|�FI��T�?U
�S�D=��%5�����m�	�E���8�&5�I����p���Bm�P����m�d{P?�нz�h�ex�r ���%*�*D {q#��n���2=/��I`��|y1D�/�0qz#�K0qˋ��'��ś��;��"d`�C��{aLI��^��� �&��5��Iq���b����T7�V��$�C�Ȓ�b �����MT�b��%��4θeC5��
���j�Y��\�_���oU���(�PrJ�sz�m�N>$�'��O쩟 3�J�G#��N�l�� H���:��6�� A��L�GP�Z(@�s�@&�УG7�<I��Z�Y��$[�б~��� �Y>{���d�Y xD|n#Nk���ݽ�%��N�j����m�p�����e��$�J��7EB7��DJ�����G
\��(��[T�-�Zc�.�-�WR%�� J��3��mbm���>�4A�ˑ
"��#�G���__���3����9�V/�a�ᾒw�|(=b]�}I=���T>�����n����$�x�D R�\�nw7���p�Ǒw�Q���|ND;>z�9t���F�\՜�Q\ ~T~Y����/h��T��������\����AO���R��O�����[�����Zh�I&�Jɿ�z����-��f�N6$b�qVG�����Vs��C��M��$|�����築�����xߗ�R���T��;:!H��{���a�ٗ����
�]CdY�}ت��m��9I��$<<�!c7t0��S�`M�"R��+�
�����Q�q�.B�b��v��jA�e�J��S=�Ʒ�P�ÃGq��Eh�ѝ�l`nqӤv�#�볍�����5ǉ:�J[S����ud�N	�&�%G?;� ̶��q�%�^һ�*�M�{xy-^���D�^7���%JaЕ��KcLfS�Q�M�.��1P�$�'� ��O���������x$(��߶��s����ɇڽh��X��;�� 9�.LO@�3�h���e��ɵ=����d��_*
���C�A�̯S۷u7��~��0���V<~������_
T��P!mHD܂R�
��b|�&��˗��U��d�9�ym�Ȳw]V$ =Z��M��YEG������>�tT{G�l��/!�D�EG��a�2�k��cVO�r'S��{�I� ?���4Tn����+[�
�9�ȴ۩"`��3'x�|��=&����GKm���@��^�@���YP׈� ֑@�!w�}5�4���BS�?G�(�#K������[{�z��i����
�bA9�ϣ���V=<*�T��$���M#!��Mʷ���RC��s�U��g����h�4K%K��qE������{^&�Z%��O�>�g*�'���~zk��C*n��&�b@9���˦��Y��0�L}�0?�kn�����뺸17c�]eG�C_�����N"`�-��H*��6Y��8i�@F�2;瑿�4$�5�g#�n�S��P�"�ѿ��8-� x���ſ?w���ۻ�9�!��R��Jée�[�{|�i݉��|�Qb��Q̇�v�2'�P����1X�����������b�
m�y8��Y����A�̹�b=*i|;! ��p�Y��\��Cʹ����k���:z"%�N� ����ة�4�򍠝6Yb�U7/:@{�w�M���LoQ|�@��hm�6s��o��Ը0í�"J�X+}j׎�`��A_���wQ"L�����4E\��j
vG�p%#w���㧞�/�r��C�	���[	�?�B �03�*��D��2���ΛGnE�����ET�ǈ<�Y.����l��7��$=U����A�#�$�'�pړW����w[���o)]G( #��w(P�Y�v�F�]mɱ�o�(ITb#qgh�������0:���'�٭�rJh϶[��~�?vRk�`򛼰,w���m��w|.�-?��;_�ܸG��+��`"�K���@��>�Y'5$ƅ�։7�uaq�	�P��G�OR���=�0�{��y��u�~n_~���Ť��e�0�m�͙�v���קVl�CR7��R���QE�J�ͣ{�����0����u��B!���'�*�