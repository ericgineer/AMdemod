��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�q����'��7�T�A&m��˴�:�u�����T5��Y�LN����]$j.Qw����F��&0�3�5�F�A�?���L�R��d��
�����8P����� NPZ8� 
�>��}Հ,Ӏ-6dvb8`�`I>;�g���:���H�f����u*��M�[��\��&���N��-Oh\k����x�SZ�)~�^�u(��=��
#�TjP�L��-�3h�(!�����Ű����?:e��s�m��oS�	��i�]TM��W�OC��yg����(�8�A?/r��>�{j�Cюv���;=,N��dVʒ�5N��D�Qc��;UI�M����,��c�l�}[@�e
r�m��<�%��P�����\��D�@o��)�����f�oAи_�㰑��������\*x�hs�ܛ�Y�e~<{@�I�-/� �
��pr⩀�{�@}�!���u�`���P/(`��&^��?�����
�^���@����IB��Q5��TKL����G��)Z[$�c�����"�I�z�]��7��+E=���qHa���Ժ��
����|\�b�K��&�v�$��Qa�Z�p%+��w��?�b\�[+��`�V��ҥ\�PWghG����aW�*�E�<����.m~�9�~�j����=\n�O*~�V�(�D/d������s$0��8�L��nUz�h�},u@.�^�h��6K�Z����M�d���3��
����㞿pb)��.�/8�^q�a�����]� ���T�gd�f��u-u����/��r��R�e	T�E��0���o�*�#��z[W�[D���E�̈́�Ǧ�Y�A\C(��sgO�Z�p��Nm�jɗ"z<:p�?ɛ	`����G�4GmC{�iBA_��s��숀�Sτ�Jf����]+�>�Lx(����ɷ�e�.蜿�9����T�sT����:��ʳ�^o:k�|�����^t��_8y���$rB`���.���ɦ��K5Њз��(j�!�x̽�ּ����Ĺ�Nb�;<O;�++ z��m��(��ӛY�b�=���.Zc5�gZ[^��5Ϊe�i҈.68�� �O@�T|"���%�v<b��t=97k�3!KG�����o������AKZ���	��O�����qC��(K��L�a��C�4�I(�''�	����y��=D�ĭS)�S�������!dLL(��99��eY<{���g�E���w�p�[[���N�rs�o)j�:Y�޴t'b6��m^�!�����{{��*�-�.vG�X���t���Sw\�#]y4 ;��r�ʢ���y'�Y �����������摉Ho�1�hv�]_��ee���lX�݄��v[��@7���N�?������X��>��W]Z�9L���O9w�''�=��t�$v��-��I������F��{}�
v_�T���\������.k�i���*��3$߭�W�G�zjw�Rb�+�ͻ�$�k��v�Gb�|`ϰen��-�]4'>�ӗ!TH�x��ϛuSx@:*�h�ۅ�3�wYy�?�|�ٮ�U�p�-(z8���a
�;TJAV�ߙp��q���~NV�q�>�t=�M:���yb��vL�x��A�� w�F8O|h��K� A�����X�e�(��2�������E�gV(�=I��@S �?ݟ���5�m֔Y�W�]+Q�&;5�����e� �_����D��{�GF������,����4�0���}�\t`��7���Gge�Pܙ�QN��J̎^���e�����QEк٫r�-%v�l}��:�\�-^���Kf�ɡ3@k;c���7E��̸�q����g���'0��k�0fm.��T��z���#�����D9!R���)�@p�D#Fx�J��Fd�ɺ�Ϥ#;(�����s��^ޤ*:ʺ+<j��G0�%_�S:\|e�&��(2������,����ܸr����o,����Z�����(V���A�!$u��->�%��ִB��v����\:U��/� ACs\j��\�uAEdg[�
i��
�)btV�oR��{Z�b����k�ŏ;���!�SF�]��p{N���@T�`[��{EAx�xy�GɅG�r���%������}�����I[���]䲩"�æ�
U�}��J��Fhy�O��S�S�"n\'��]E��I�C?�yW(E�!�}�QG!!b櫩"2�4��E�sӒ��(�))�.tۥ��]���;��Ӌ.��W~U Ej|l�/T�,wׇKG4��S��b��S�?�?¾�C�"r�D�H�	*�.Oj8����ɪ���q���I��v�v\���88R�U%/��[9#���"�����jgы*Fbrnv�����S��^K�9(_M��$��%��δ'8����{`�7���ئ��:�5��29�;|��^o�z�v"��`�䔸��P��O_j@��nz7Q�D�{����zF|E�3�����2.^Mx\r���x���>V�����^����	M�{��I�%$�5��6j�t-�(tv�K�F0_�SVN�b� P'`��Z�O2ơ����1�5��R�RNm�)G�Mmp������sב+/� �aL������<��ą��n6������@��q:�������.�S��n�2���a�������X���p=��K��;-7�9V/#_�p�ۂg/S3��ymRܖ�CMD����VN����<�sO<ZŜQm��ޅ�OI~�˨q��jS�<��nG�t�S�'7�w�w�M}�K��-Ym��L��h�"��F�����1��+�8{���0�U�;'L��ޯ�X`m]\�QD����*��(Ǆ��{�_� d�gRp��+q�����ql�R�t�2��:$b���G��W (a��Ӛ��~�!���>��48,�v�B�Cldy���-���۲~0K����A�Q�6���f���G�{����k6���&�j��gJ�vlv<�X0M�{���׃���n�+�2���;�̻��h����|����eC��y#�eቄ�%qY�Z�?�n�G4L-1�Z+�P��r��K��Ű�v�K���[���:�Tx�Л��`7ԑ#;R'-g��ȭ�@"�/���H�ݤr8�[���m6���]y��5?c�:Ȯ<t��p�_uQȩ_)^#Ů�¾��g���y�&NhɽYg��I4�PVp1�8ChP�>��٢��Y��5A�e�������\n�h�� R�����	^�X
ܡ��⮤Cnst��B�(�\�Ъ7���#p2��wG.E��P��H{�R�γ�]pbSw�~�Ya;�6H�GC��֋�%�R���Mw6���\�6������"��<�Ċ�T���H�,Cn6�P�Jf��7A1���ئi½��(�ׯ����ג����n�'�Ć'3`���4��5��-k�JV�}�?�3W�4�Q��}�:���R��gι�3S,@K�����N��7�_�᷸Z�[a��e�zVJ"�		��ʖ�g�Z��U;cA���l�\�8�r l����+c�쿮����CƂ)e�w�Ks��e ��>���K�b���#&S`4# ��J��[�iiQ��5Y�]mޥ�d��]ܝS^� 6�t�m�J�y�#����{2�����U�kL���":�������[Ji'e�ڪ-�1�������m�L�]
��Z=xף�,�W��C$�8�{�Rbک8)�!y=�/�?vѲӿt��Yx�u���  c��'�sCv���ju��͹l굜�ѢpCW
�_H(;���ˏ��L߸�u3>���u3�M[=�5!�N���W�G�������x\j�mѵ͵v�����g!��c��>��c���d�S��x"�~CtG/�W=��!@g{�H�܅�e;���I�M5�x�)�V�N������"ҹ�C��]W�� cR\w1@}���Y�z��#�y����-���������xe7��'YU	��ؓ��҄FE�\��_蠟po��5�7�Bɕ��r�� �.\�
3G8+Zo6�m������������O(��[=K7Dd��w#��/[�u�;'!k�6�h��lg�9����|��Vܤ%)����b��J}{�j�ۄM��yҩ���y����رe��ق�� ��!x���s%��z^�m��R�O}*u�4>�X���X5O+@��m�cj��U��
|
��Ȱ�a�:�F�~�N��}:�jb�3r��k�/��e�9��ߑ<���2�߫\�1C���׵I�l��g~$�h�P�>�/;��D��