��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�O�5t�"�/�V#�bnQE{C��P�oHȥ��S㌰��'�@���:K���J�7&V�T����F]X�J�ʨ(��̰͑ާ���bރU����B/,d�{X�F_�@�v�k�7S�x1�=�2�T�ޡC�� 9$<3�W0Q���a�.+:��JK&&N�O�6w.DᕻW{wG#�nI��1��҇��P���� ��~��y�i�g�`����7�E\c	g2m���k<��� 	�Sj2 \�F\l�]:�/�u!hd���ڬ��'�q���bVi���c�r���P�c��%��º��(�'}�2^��6Հ��MVNV�
-xTNI�h���ŧO~c��	���P0z'r�r�����O]h`�"~�^Eݺ+��.I	���f����7���.7���\�N�T4sy��C�Nq�O]�H�>�l�􈯣��spx��3��Dq������k6=�|�@��ܦ�ui���v�s}[ߖ$�gY����c�\��Q<e��I��|��xk�;b��Cg���q�ZW�t��0�Gӷ��yn�;(�=Y�����sV�Y�o��3���.,�I��#��֦��1�k
r}Ό����^�!��?l��Q[�D���|R���A>ς'�L���Ŋ��ȼ�����f��"�-���x��=�H�I�ZC	P8j?0o�!Y¯��J;Fr/Ð���ٮ����jPkh�G�
�*��v�j}i;w��^�V���*�b�aB�ʸ�N%��X�24��*�}l!�-�_X���Bۅ�/m�/{����_�4�A���}�Ì|�V��v����p��(���##mF�����c�&�7�hI�e�?�᪒1��B���f���>n��Р���G�Fض�-$�>J���)�%.XG�oJ�p3Ll�(�rӍ�S'�N�F�GB�������=�V[�$2�#~D���Ɂ�l�u4z�@��@�;�+�8�i����QKQ�E�W�kRث}�]%�m�aP��wƋ�6�˹�9�'���� ����ȴ�P�8���-=IY� $.�o\J{C����s���*f �\$�pu(�{ޓD�I�&�w[��5;J�J������3s�&��_jN��1����N5��JyZ��|�)�[B�S�Lrif]ٰ�b7���u[�9�w�$H�~FT��5�Z�W_ � CNhk��v��kS��$}fۊ��u-�	ͺ�2v�eW��V���b��e�J�]?��,��Z� r��B�ꭲ���,ev.^]i����VAK�(p���yo�������w}�,O��&�Bɾ�Cu٦〹���'���ř�޳�2!nu��Q}�+\5Lz��_��(���dqi�PNo
1�׮�a~���VXLg����+�c햩�pb��m��w�%��bx�\�+�S���#""�%(Nm)A�Z���j��$�f?�L�91ȩ|�H�L4Tc�H�W~;���*�2g+���GN��d�+dp
���p}���j:7��N����_�ܾ�����Ϣ ~\u�x ���x͑�$��#H3!6�c��mL*�Q!���!ұ��z��&�I!u�i�9�*!?�ηJ�G���5�K������>�c����Zz������Z�#`�7���ed�uyW8���a�M��9.V������LD�Ve�&�ʏ`�x-�V��}u��G+R �Ui��(��ǣ� 1��7��4<����	��xHN0s2f��C�k��ΑR���U�o���U�Nb���K��.]!��i��>zE�<�MN����2��9�+9����;����I)��:�������1�c6��V�n���s_6�P5��F}�|��� ��N�]�X�X��S#t�83$�{Z/)W��":�4�R�u���M9�r�Rգq_vL�ޭ{��>�QwĮ�aQ
X���]����`�i�$��Y��m-^�����N6�C�8r*KU� �a@S���!0���h��Ғ��SЌf�Wq��2�!v�n���d��a�,y�.�tqϽ��Wt���D��YY{{��]��� !����n�Ŗ� �Ál��5��7E�ڱS	�ݩ�H�(��;L�T�`b��:NN�`�VW�1v������^���M���f7J=+i�Kya嘹/~��yz0I�;^NC��1A�B�Q\P�~��^��}<�͙�c g�����fп��;g%

���3r�b�K��ؓ�`Ҳ�Z5 դ?��[&��9ڶ�9N\�`���y�:<.��\x,��\�[�ñ3�4�C��?$`cnU�B.����`m�<� h��F�32�G��W���
IŠ�\��ۭ�(��*�ZS�-W>��w�o���!��%������T!j�q��m�8ʺU/Y;E�-0�[4��:�ˢ�1��muu¹�V���0$�Fri�����YFWAF���+�z�����:3{ka�v���2��yj�!�75ko�8Smr� ��g%�������1�T[_ O��c.[tS���*�#��<�&���Gڑ�Ӝy�*����d<�W��.1t�����t�t�HD>�|v�u�����ص�3 ���q�Q�.O
)�"9�E�MN�w��k;�}I��A(�����cc7GM�BY���� ��<����Fw)8E���5�o�&M�)h���ERZR��6cX���,H�.&���O�$���l�@�-=�^�>�����U�N�:�i��m���R>_��\j���o�n��G
b�ԥW�ݦ��}�����z�i��"�� �>ɡ�u�vY>�#������~-�}���!�� J�����p��O ��7�/�;硋0VW됦�V��?��,���ir�{[���-���t��p�`�	�k�v�s1�����W��^#6��񜕓ɿ}mH����Nxi��n�q� ��@���M_���
'�X�ɋ�W���ǘ����,�S���2g��[��Ӎ��ʻ����Y��=����yػT�0.g|<�ߛ"�(�Y����,���)y(Җ��՝Vɡݱ�j�Y��6�v�]�w��J�4��o���3O@�I��w*=w0;+��7ؕ���\֢�N�A���G���q��y� ̑a�h@�I�Y��[@C�z_�J���&��������%f�]9�H[g��?��A��k��\~Er�B���z�9<��zǧ�������6�����
9��f'9�����R���p�j�К�<������VѰc���.�ّ})�|a�M�ݭ���7���ä����[��_=ѻW}G�vS�����Xܝ����rB-	-��`g:?��y ��A�d�~~�GG�J�a�>�%lU%*T���;4c��\/r�f��=$��^t̡��^u
�V(���s�~��ޟv;D(�Ά��:" l��&��{$i��i��v�n���3G���ɿ*a�6�Ȉd� ��7�)�ܚ9�bʰ��V�N�v��򈘢cb�@ڡ�wYb{��d�)%���Z�(/ _8�ݖ�J������kMo;�:�ө��H�'��/�'H�c�Y3w�B8�{�K�B�-H��!�L��+:�ԔJ����i�����V��v^��,Fha�v3���Ҍ�"羫�4q&��oU(9�F$�X!��t#�3R'����V� �y���8�D��|��-hT��o9l�.���i�=Q�[�t��Ms��u�1��>���Gf���E����r�G�v)�h
�5[��MJ��+oo�;[x�y��?��ܔʦn�_��W�a���['�R�waEɩ����	�����mߴ�Ͽ6H�� q `��U]d�SC���(|]����撴�����Ev+K�/����rl�9����k:��hk�Y��Wi����rcY]?�#TK�܈�C�0�e��m-�2�"S�@-��WPM�=��?i��DPAtG�p���3�@/��z����me��6`s*	���EJ����+ Iђ̧�J"�(��#�_l6��K*�D$����q�;�n>Sy���[I5
Crz�g�rf/ZI(��n��W�LT�D��JUb��6�h���Qo��9��U�XW��0J�'RS5Ju.�/+�V��=���V!o�?w�-��)x[y�Z��#V{f�Y�r6R����H�s��e�'���Չ�w�W�y�uH�:,'�Vf��%|�3wcv���r" :R�i��@��6f��zf~�,��5���3�� �L;xlz�Se�ClHY�~.OޖfZAG�R�~�$�s���SNZʉ���	�n.e�4�"^��3P��;�R��(N�q|oơ]��x�e.�G�!����~<������s����w�	����S"OA�mv�?S��S�7�HKgƱn��WI�o	+��mЄ�&'��陼�j��i躾�M�����oa�J�0O�cUZӊ�.R9���<L8sm�s$�07c_g]����mz #��3\`�ǸBi��&R���J/lD��n>�j˂��1�:C�#���B��I�O`�e4�Kq\�:q[��D���i��]C�Q��\.Q$��`=�DE�4o���#y�E�P���H9��<Y8��!�7{��1�4�G"Gk����8�k�&�hN��,.}|3%H'�YZ�y�䳨�^	ֿ�"kq��>�#�&ݢ<�v�M@�,�Q�uC��g����Rӓi�k{@�]�� �xQ�%��ه��_KH`b�i�A��^��`[�%9æu��z�k��p�F�!zr�{ޗMޡ

H@�QT�]鿜b�`�T�_ƈ$�*��'���pMs3��?����GSt��̐�}x��3uR�q���!�J�.˝jJeEuoa�3m=7M�+�v��&(�����/~���J���-!C�ƥ�:< ��h��l�lg�G��_�L@~�/��&]�W�ܜY�P䟮�#�K{�.=��8����U�l��&������梖��:H�Nw���<_���I��-�%�3i�ᇂ-�a�Pi�9��=�D�D�A��D��F��Vpcu0ט7����r����۳�JF4� gn� l��㱐��ýb둴�P�l�������z�˭О�W�TJ��¼up���n{�\�3�x���~��R��R(��"����.��{p�� EHaf�	o1��p��2)�n�������N<;�N���ϩ_�k��~�|���j�fg`1x���JV�EM�?���M�gYZ3��j�\��?�w�f� 8�'[6T�Ӈ98�4՝#q7����X��6LR�TRdN���X!�l�����B�@��K�f�Y��ٜb�'z���#L�����ܗj���Ƴ��}N2��-�.�Ǡ�Y�]̗�LG�,*�JP��K0���R+x���Hv�i��5�L�j��B�)biD�⪕����=�*-g�j=2�����L����ˁ�}Q��<A����D�_�t�ZDX��Uu :QKI�H((
@$���i�S�+�6f�Фl�7ݰ��bv*�*�CM��3�UBx�-����\Q�n��jk��h���)(�L���Y�Q[D���e�P���4KF�{���������NN��Ou�
q�M	�@t&H��ۇ�+�nF�&A#���e�tP�kZU�[�x4ӹ	B��7���}�f�b��Ҥ3'V�
F�^�	0N��	*�%,׶��w�0�OR�b����,���7�0�'w#�a��Sբ������EɆu�cӽ��)�t�l	�8F���m��:|����V���/	B��]ۻq>ה��ǒ"��e�����L`BLؤ(V��1�m�~��=$be�v/>/�~��˂�[ύd4iԫࡷ@=ؙ��)̛�G}����{�� �������߰��]ϜT� �F���7����3 C\;�i�<3e�$ѩˬ����t2"0���#��%v�/��~�j����b��s^�E���3���1���П�2)kP�ky!9yϖ���z(r��u�}H>��4��\����{�K���>���9�T��x��HC��ud�ܿ�'��ůW��� �t����@AS�C�/sgV��Q�d�� KU���^C��3�C>���(������Q*��� !Ey� �5f��^լ���]j���д������nc5����@��� 
�ik����� $��2��ĎL=��P�t��\�itf�}��L"կ�X�m�4�Ǭ��A#�㭤�D4��!�/�e6��y;k7���yq$��m�=�	f�R\��2�����]D9�{��%E��x���|Ec�b��G�H�s?�f�OrZK=�1�$]vc�*%���1�� ��M��,�A��=q��X;�@'���<��XAQ節d�-�����{ H��󕈁��T��d���w�s���l�mQ��$�L<��v�$q�	c���<Zfr�]�,	7��NEx��'4�#� {6)�:+8K���H�t _���z�w�� Ү4N�,�6��{����7f�/�~'��޹��캘m��r",�I-VJI�,ugo�0��/��Ê('�J�cJ�졐D��(d&��r`Қ&/W�	5^����ye���*J8��	�ŞɃ�>_�|�w���H�el��K��2��k��u+E{�O0%�%���h:�P1���ÔjN�-�� #@�=�Vk�[��Ě(������ϭ́L��υ�˒�q~r���zZ�2�h�����鉠�;t�:
��jZ�E�
3m暔�W��6@��I=	hЧrI6�΋bU�s(Fq�"��ʍ��%E]�x�)��:W���75:�8*y��w�j�Yk�ކ����Z����GS�O�K� �]�.����o]���ouG�CĤ��`�\�L�IO6�u�X#_��/L�?��6�U�¼=�y�Q�f�,��t����΋�R�v���W}]��0Qx���Y^*,jo�M\���ׅ{�_X����z�.��a	�S�(S��h�6�2;�2�2�Wj��_aZ��?u�i=�&��	�OM�rٻ1d�ʾ�4��B�j.]��WG�,���맾�\�ߵ�N�:����ca�5$p"Ҥ��y�	�D:1	r���|�g�ء>�|'�i�!�RW��������[�/���J�j�N�t�*{"�����S�48�]�����V�� �\h�?�Г�+0����C�<���Ft��٠��7�e��A����&,N��7���ˮXM��:ޭ�k����:u
q�Ŭ��Pb��*��(�I����J��Z!�^���S�´I��ܭc��n��wX���a?����-��(��L|z͚A!��m����,P�(�F�Z��kYH����~��7:x_�@�Y:�%er���D��Q�Q_�g�\���ֺ�p��#+ 46��A�{�Yi�3E�}�X<Ӫ)�7�C��ҖC���E�A�!��=����������Ȃ��S9�W�-���yiT�G�@Ʋ*/d�*�� ��@Y�y>p�>�^�*�o�Y����&��F7{i���$�΍O�=����YBK:�Kj�E�Vɔ`~�����	�}��(�B&u�S�^�[��l�6�@�I����h�X�W��gY�<�W��>�{���h�x8�u�O��P�<�UO�/��c.N��׃mLU����/�?��j�1B�����\Ĥ�y�Y��L~'cP�K&�"���;����!�gQ�DU�t��H̻��)�]�sԸ�����I�ԏq�0�ux���Nr�; �@W���%lTw�V`�֔v.�+��ͭ;Emxj.�5K�ͭ�id&]6�sh�V���w0? ���Pa�8���7߸q<g�ც� nn�]��M�XV6�V#U���1�ԸbUo��ϗ����{Ɛ��Y�lq3:
�0d��N�@٭;\�%�3
k�߱^c�VK�ag�c�Ñ5�M*�g0� �m�P���"�eE�<<CyY3�������i�G-��if�k�I�P�`T4Ɔ;C�n�ͱ=��9�N�욿�_�-�~����iw,D�I����/f��F�D�A����XU�0!�?���n�'�A�
j�ƿӝ��\��~!E� �v� ����D�5o���{|m���i���<$Ygs�u��+ �%��❕�6�����ڨ5L�d��e4c�Q��R�!�r�B����#���*v�������J�Ւm�M]����P�5:��4����Ì����`����x ������H�x�������Ks]�&;%����ؔ��©���j|u�}V���$�T�ّ���;�cy+����8�#o�
?Õ ����\���/������=����Q⡘&�'=�D^YN�cG��ɽ7/���r<V:4�"��[pw���5w�L�.W��d�'��;�Z�����-�Yg�=~)P�>Js �}�~��M�C_AC�������9g���1bZ�]���6D{�T$U:u��A�#��a?��r����Z���F��/B�n�����J��	�d^���~�c��G�S�j��\�&D�b�[a���w.��ot�����/$�?�Ďq_f\p-�#M-k�i�2$��G�V[�`�Jh�q}R�yR̊�����	8�;F���3�/�wH��c|�"̜Bn��ak;�\O�� �Ê!��;�Թ�y�g�N@�6,+��v��f�9|�w�x$xJTA]����� 2�^��g�����gi�^�/�ϩ�sD3KBtQp5��Ȃ��#���H���@���9�!�u|�Pm;�����/�d٧\�R8т�=x@�x���-I�B8هH ��i��x��4	��Wv�B�3���K����~
�ᢦ,��T�`�T��ʘ���CU�������Q�+Xߧ�$4O�j�@ ��*��\�!���1�.�@�{B"�ڢ��h�<ͱ�����v#`��ZV��_�M��SFK� �Q�9���nI�%o����A�EbM8��2�A��)�J��E�ۋt$�n��o=A�r��2r�2�iT����$1�/w�]:^O6c�����{��+"�>;Y����ƗK�&�h���
��ㆻZ=�VSX�p}r
��\Xpe8�1�'�t|$#����yV�Q5��g��	?��q�曹L�
-q�V��E���SQ�s����b�W�[9���Vk����ǯ�J}��I>4A!~�4����F|<:n����(BA��w�l㾦��d>�����?r��vQ�=�1a.*v��2R����`v���@d��-L����HY�y�<�;� ����@��U���d�浹<�,�P��'�&�k����-)U�~�
1Da��o͢7����K��wD]в������cs}Vn��g�9�|P�� �0�*Q�B����5qO"�Ȕ����\��vЯ��B����&9{?=_9x�U������P��Y'
"�Fܪ;[-��g���)�a��m9Z�V�OtἼÛ"���o��ԓ�+��煾�sW��"��\ugJ �!���Q;˲�4=�6���U��=��Y��E��O(�ի�&Ɓ�I�%�vJ�rݹ'	����rʠ�"����	1<: S3{#!�Z�z3��	}�����t���y1��9r��i4L:�k�(�тBL��#�f���b��RD�}���Q#�h� ��hJ�{��Jڔ�i4�-�˭��Ď��n�Ԉ���t�x|fӉK��p!�6�u����ǔvʒ^�8�8tϫey&Q.����(�R���鷵��5�Z�����LA'��'4�Ǽ,�#vҿ.sm��X�1�G2��J���,���)5�����D�⇏D�91�p���h�^g�ܗ:�(��;����XBI���c�D�<hr�� 1k3AĖ �3���&�W�1j�3������z�	v�d��`I�����A�(a��'D����%ʭ��=y�M���bp�ipUM��Z@�~	H�V�$(Qg��47��W���gx�}��C�AT,ۘM�A�U&C�'�F�D+�[��?2���pl�b��D}Ϛ���7���_�Qy��Lb6f��1�� �Y�?�4̗`�t���6D:����ht1�(#�8�L���S�u	�Sk�A�Np̂r���=%#q4�*M�s���X5�`o� �eN%�B�;���p̈�J�z�>j���+S�b��5r'c��3tA�ӈs#�J�
p:fU��j7	����8�Ŀ`՗o �f���T��XpT~�j-�m�b�e ���S'��E��R7=��.Ȝݫ��f8O���˿P;�ՌC�/f�x;�w�O�������7��=���Ϸ!�� 7�b��k9�~��г5�~:�!sl5��h��!N7��D��V��/�B�u�S%���'�h����6�yOk�Hh�l/�Ӹ�p''���D8��Z�q�v������	��d�nEn&�O��X�As�)�B
Dy���?�ǫs�X�uV��ݼj8?(+��,I2d��ޑ`7z�s�M�+:�:�y��3�	���i��L�!��<���B����iت�ן脊!s�V�/�j�/%r��E2���Cs]ve+,�}db�.ky��-��eE^c�j<��gF��9�	���T�.z���l�?�M�,G5R��r���̧��ڵ�;�9��콢z���=P݅�%� �����M{G�Qs_�QAQ {���������Pa~h�Ѻ5vv��%d�N���M��@c��7��'���D~A�V-���ºP�n>G�T��nV���6mϜsv{$ϿPaP��ʪ�$�fd���N�4}5;G$^�/�d�'賂��Cv&�ۚh-��59s�c�9����lF�[�qiB �.��[�KJ�ē�B�b�o!�Q�!J�d�n��tz���c��w���I�����R&�p���)�_����Te�XNML(����+4���E`v	�����ȵ����������g��Wrp��(����ʊ|fxN���p]�������+/��%ͣk�o�ʘr������dfə!3�����@�M�G}��ץ��핱�3�2�vr>�HhU]%u�v������ud��4��:[��	p7������J|�d'��q�*��1�`A��aܨ�B�a�hK���X~S�.��X�z�;�9������(��yl���6Ah�}*�`a�Vx�u�O��\�Ȫ.�a��d}x�BEwH�����cn�=R��V.͛�,r�G-��|P�
�m�{l�p����l��k�{I��|3��*�9~�.[���~Е��I�S���#Ƞ��*�N�݂��Q��c��s�OR�`ar3�hq~�aQ��~�廨��C&?���d��o�d���5�- v�?4k�;�?��Y�Y���5�!���y"�[�`d�sE���.�I���/z�o.�%�[y��\_��>#��%(?գYE8<�VO�N�����[����1W2Иs���?���ژ��<�(�,�g����O�F�6%���k�=��@�NG�@u��#V0^M��1j�-�.}8 ]��������݅r,}T�\��;���\��v��8��5�@e��>�oo��M&�K��9JŮ��M	��CL:��
�y938�s���N���?�ɏ�oI��� R��������B�t2^�����T��n�F�+u�]5!�iI�~�Я�2y�8��1M?�XCL �����H��v�/ۺ��V#�\�����-(��|㴸�U�_}U�P����|�Kx$%���D�7:R�2UE��ΤLa��0c����X�wȨ^�#����DsJ��kT@��E�I�a��p*?�~��k4�b!�K�b��CX9�k{/
�P�@\71�Zm啗�Q������&�����&U>֌ռ�@\�Q�p*�ًX�E�oiN	-���
���'Y+��i[��&�e�~]ETZy�1��L�P����1���Jh��l�m(��:^G��ʶ��B:l��A�)��;ǩnr�j����5������=�l.��*�|�~8&�t�@���܌�������ɺm�~��\Ì�Y!�/ĩz�ok�trw��i��^r�����vz-k�
H��[K\ #W�'���au��4	�5S���h�(�vM���_����:��#F�)v}9y�G�wpCP?<	;}]s��!�}F���o��6V����xo��ڼ�e��<�{7Z�L��f�Y�ƸI�Q�7w�N�]ɳh=�G3�ϯJTV��8����!���?�8M�����֏ם�
����	��A�3���4l���#�����?ÉQ��'�%qh$��R��4WA�4G]&�U. ��V��2�����y ���'ճ�| f���$Ȫ���1rV���?a��ту�c���N��WFST+6l�|�_9��2Տ:͛�T!���GD��TC�ζ�uI6���`q�>��
�)HL�bQ�]ن����@��K���U7�d0c��{̰#�:^V���� �m����*�/��˾�\��&�*
g{�`�������������h/I9��鮖÷T�,��j�;�/�hE0���_WZ����:RW�����p\?Fw�3�A@��QJư�`� �Rn�;ʖ	6?�K�7�]H��ݽH֚)8�C����Q�c��Di,�� �IH�UnO�� d�����R����X��P�j@��i%=���q���7X$��}G�q���>tvC��Q���#F�ʙ^�#���I�m<<�ݞxD��1 �E�PH`�1H��N�Y��D����1��&��)�K�F�SC%�v���	K�-���ÿ�P�ǿ��t9W�=T1��2�H	�O
5��T�`�1��Z�4r��d��sl��V�Y�����v9�[g���sm�bp^��f�P:�T�xR�.�oOq�;)ꔙJ�*������^(yfi��m�-�HH:���VsP�-�D5N�1-�=���VB�H�� L6Kd	��D4\AG��ę�8o�Z�?%{V�V87ؔ�����Ph���ޫ&�%蓺C!��b(Q!�,��)X��3�Lb	���Y�Tmk��(Ƽs������̠!�r>��[m}Z���a� �%���#Q/�d�7m�����ZHBy�/d�@�'��S�P���gm��W�8Kb~�8
6~�b�|&����3X���@���2o�&@-�B�����*/��喬�����+��A(�g����w� ��L,
�!�)ٓX���効#�Z�����W��)������j�9���$4���Yv�ǵ�6&7C�l!�r�a�w�'[ܽ=(͇�lʛ$���7쏊����hPH$dg�
�>X�:W�C�q���a��䏵w�n�89�߹��Ķ��qH\� �;Wؙ]��}�f,��8�p���/=����a���aι�m��W�e�n�7����.q�<�^:ө�g 5�Ï��É_�U|z���f���cu�s�~�K����}�a�7|k?&�"m�#������¥?9K�Z]`Pw)Ro�7;m��;(&�tuǮ��,�3�*�����Y3k�g����9������p��"��i��=��&9�(4��{�F�Qn��q+��푲���A��~�����5<�b(Y�b���Z�I��x�S@#��s�|� �uR����!Μ]i%�J���}v�R� Z��@T(��<�N]À�4(����@̼���p#ݢ��u[ܛ�uCj�A�r!%k.��s��2@]�O�'�KO�s��|���WH��fD�⸮��ב�=qx����c���A��ů��s&��q��'nx}�:S���l+�T��C� �@�y��{��|Χ3�)�O��Y�堁�F�P�$܊�<���[}���#�Q�Vš��>ot�\�8�]Ȣ���Q��X=$"�����`:��