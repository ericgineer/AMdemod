��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��Mg9��X����6���
;gKd��Z{ferbwN�m��P5%�a9�/;�ۜlڿ�I0(��Z삥��*T;��3���*Hč�kOg��L.;v�ȫWr�_d!��H�0�/���d���Z$�OV���hà
�3���w�� ���;�	_�Ϲ�����\䌕+����0�l�HϿܠm?�Q��\�ՙ��o�Пoʻk����w�=P�=�C_��OF���S#v�8���#��J�|�H:�@�U[_��}^sK^���g��|�7��x/��_��N���1��6� 恲@�)�.� K�̟�҆H7�;8�w`����0P��8�G`5�Y|fd&Y����e�#B_�PxIkof>����y����뎒F@�}����������$ "$y*#�F����$4���ſ��Jqё�������ŶK��/��ʤ�����/�E�i^��L�AH��M���<�	��=�ր�_N�d:�7��U��D�-Z���y��įiZ�ӳ�45n�K@�+����S0N���:7�o8nܶ�NB2�֤a�ӈ�����`�a�uR��'-�di�Q��{Ǥ�B6����h'E@��ZUJq~T:��ăiZ�. �⸢��i��h/D�����Α+ŝw�$�q�P�M�C�Sݶ��/r-k�{hn�#�����S���%*��s���&�踘C��4~P^��C�8>�]�s��^F|O]�s.��͚�	.,�
-��+\�V9Y4�r6
������l�B��˓Kj,z~w�81��R�����@��73!�9���k|�/��=0}a���Ȁ�L��������2ک9	�m"&�j5���%�ʭ��CKC�M1P+��>hZx����Z� ��sw�jV/�{�K�w�����q{�:I�a#�ĥ��S�`���3NWhNNC�]�����PU�	�0�Y�z�-�M���ΠO%a-�?T�6iO��	�g2h0`:�^mT��17����T��;��ϡCq~�}���1mb9P�ȟ��.@��,��l*�s9�N��g�����h����frt�_�f>��b}��E�J,�;=T82\�'�ޫrU��Ǒ84���1��=�~$+�����B!�P�yז{�:�Y���|B�>�%�5�ஏ�Y��a8\9�7W�ғ�G4D�-���S�|F�Y=��|7����c�X��aA�E��Bmik��0c��$Y=#q��w_vf�K��h��w%�t�LF9&<J]�m
edHărd�bI��'o�	 g^��u��#�ڿQ0)8ʥ�2((���9j QB��k=d/ׁ��	[ux��c��^��\c2h~@N�,�N�fd8�+mB�w�|�i��;�I������G\( �x8��JV��-�9�m�9O"��W��h�
�Zԃ�k���"���[ j��G���cgS��fy��*K�{��"rFH����th�ǃ�p�^�Q�I����i��c�`t�[�0���NZ���v@,^�αm-��k�y?�y�M�HǢS�a�
�<�g*�=�^(�1�!sE�\�vb�&�`�z�KH᡺F[�9j,�	�[Jf�
�~ʑ�{t v��>%�A(5@T�'���c��3_�XQ�Ϯʤ�e�^oʹ�e���ShE�=x��Cm��I��Hs3÷H��A9��d�z��;�$;*�iAkW�1/�օ!��o,Ы�^�$ʘ�L���4o�+�Yvz-��&Z�ƴ@5m�ϧ)9I
p��N���k�5�u��V�. ����<`� }aT�Vk�cg��M3���Aj����ő�d�sŢ+��_N5֢N�>��,ijà�{�tA��l0�2��,)V�ȕ6��Hm��6ۨ�o,>҈Bֈ��j��
��?���C�O)��^CI����'�#�A�ݱH�MH�.?�Lȟ0&���:)��G	����[Q��2��Qk=�I����y݈�T-�4�I\�o��8��1n���R�I�4H���Ff���-MX�Z�$��4J�(�{y��5;��U�]��P`U{4Ӝ�	��6�)�e��в����#���Us`�蝇єwJ�h��)�l�Lv�Ħ$~l9��냁��V2>��ݬ��)1	����_��?'8E����KU|cs�~bMِ�T�U�4}�����5���R��r����tk��b�}>@�`
��9�-����	5
u���-�e(S�d<��8,��A�s�:DG��"�,�I	WU�k�����:���E��d67ꓣ�:��2o���6�v@bH����
�2�
�����v��e	��~��%���oƔ��n����۔��� 1)@a�u��s�D=�J|����>֧|W#��8��p�KW��@��v$�)m���Q!��{W�x?��9�b�,O�O��}���]"3Ǭ�y�/,z�m��u\��J�n���9��W�����ӛ�V��v�0�GQ&/���/K�����0�d1 �F���Uȝ������O�ݔyھ�U&�c@��B�L����=Y�0'��T��]@�"���-�ğp#~�|ٓ�q�:CƓKk�ۇ*f޴3�E�8�{��ڙ���w��Q>��j'�~�^m�l\IcVTU[C�ǳ�Q��4۞&sԪޟq��ħ�c$e>������q|�E��o�oZ��YMa ��<2��ͧ�@�<�pE�g;G�t��D�0�%��ΎH�J)��;��R��+B`��dH���1��Q��$�8$����-���mG9�/vk��y�u��(�]�4�����LNV����cp�B�[M֞�4B@(GD�?	Q+P%{_�����I�����o�
�H�Mn�o��Q�����,���Q]S��c�K$.��mp1�+i킟cET��>��S ��/��KQ�Al�P �����U��5{�o�j����l��u%*�J&���Wh43������k��R��3��-D���� s���w���Օ�?|¬/t����O��I��Jg�����a#?����v�C�y��xd�4]�凝aiS�����y=<t�ԣ�x��<����}����U��S�B�3k;���'3`��y��ӘC�;Ӵu�mu�]	�E�+��f���"��q�l�P���^�._�=)Ɵ�X#���JS��A�� =#����R��a�Ҧ� 3a�%@c� R�S��@����b��/�"sa��_�<<U�kMK�=,Y=`�i0q�E�d��B��|�͐�t�2�٧�#�����t��P�8������l�I�U������<N�Қ��C��vv� F�BX����>T=О>Iq�6~��'"nH���9���\5��s�~"%{�Y�h����Cަ��
� �����{�ʆ[[r3��F(J��ȶLE/�p}��A���"r���y51rS&j~c��9t�(��)�p��B�8Ԧ�
5��Fó��c�$�JY�!��`�$�#�sʉ�Y*&�}�E�U9��T�|�ƤhA(�C���OY"��q�uRZ�OI;F�l
)�Ct��2�O!�O��|�z%�-�/?��ݩ��J��[&�B봿�g'����V��=��������fY�mw��A^�)��8�|V
��0����׿�3�e�}�v��;�._<r��,�6� 	9��"^�r̨��?��Y��NVXZU5&����.�!9��)J]�%�\YT�L��f�O�3E��3ZG�p�0�w������U�w�&E��ꗩ!
��%o��P�ݎL��NLG����e\��o|r��hrw���!����!Zr�>P�&Ԧ�9§o㡯�Gŋ�����"�v���(�疛Ⱦv<@3w�VA�I�,�����s����;�[�Bk��Ŗ9��oWIwM��7(X�F����{���X�!����FL���F�{T,�KQ�Bͽ��]B�-ڗ*jѵe��w�E��.��A����%)�ie6=M�t�m6�:'ns�4zgֶ��cV�P\Pd]�ޅ树\>�-G�̀�9CC�zTG�:�w�r�&�1|0Td[.���k"��O\�u1���9*F��������F�^���1*�d1	Dw�\sBo��3��,N����%�kš�L�l�B��t	ַ�ው6���Sm�+�"��*T���2H�붻v�]A�~�I�i`ZI2+�h���7���{��D��fsz;�l�ƿ������H9�A���]���1*96���+��zf�>ħ	 Q�-�(�P��}�B$B�<���fW�`�ǌo��?*]��SZ
���=�I��Ҷ��O�<��!7s�W�r}�V���a��pzӍ����R�ii�2�1�\t��w����>�L`ʎ�7h��*�#-o8�W)�M9 n�`��A[�8B����5�ˁ�٦Fr��~(E�����P����i8�?��p���S�H���k�]^�9�f��#v��1F�t�&~)�����s�%�@_Z��"��jyd�Z��f��>L��_f+�&��� ���C�q�il�����c��}��e����������*�X�DVG9Ģ�����%�U�����fq�ו�/-�a`��Ԗ!O��sr�4{r�f�p�B�w\]���?�e�E��Υt)�7	��*_p�F<���(�dڗ"�2	BXg\e��"���m7�=�>-�'l4�O!�-Q��z)���; ;�z��Dn���~�&�Q�( �"�*Z�3X��Ʒ�Z�,�@\�P�S5��g��g`��Gt��?r�j�M�fi~�t�WO���U������c�=�˻,,CZ�3�g{�W"��?��a�|'2�#����kPph�k0p�!E��,ޅ���*Lz3�C�M��)�% 膄����.mEa-�a�*I�Ғ4g�ߤ��_����������zĒ�$t(ZT�ފ���	ܕ��M��)���w��D����L:�������6?���f�𲍶U��)
��{v�t�z��!*z�a�msp��x��fd6L��N�:�W�"�0BD��^�<�� �K���\k�Sƻ������;�x��qQ��L�rnIw�|N��]0~4D�Ԃ�¢#��������ƒ��:�nE��ju!��p����O�R­Y6�h�FzF9�������;y���D�����*ԣ�p�w߀��m�Z�3ᔿL4�3�%�T#1>Q�E:��|r/�
ASB�5�*=@k�j���/���;�?C�1��7�D�A,A�z�<�aqͦ)���,D��w{��S�?�O�:tJ���m`��P�nl��󾃑��~ےW���b�f�j��M��LȞ���D��`D��8a�V�y��ʞ2�e�u(\�ǀ��7�;�"�ʅ�)�3���gy|8�}���BAǄ0=l�����.�c�w���ˤ�i_®|��3,��@�8��[n���C��L�1=�uX3����t�PY�!}č�L9��2��~@>{`Hq�/,F��c.��=�]�R�$v6Z���K�Ǹ<���^�'E��D��َ<&���w���R�8p�gU��r��A�!GO^����7?}���fރ�td����=�r����cTN��c=e!�A:t���з�7M��>��r��`SG5�nPDѬ���K���/0�&�G�UYvY���-W��2�i��50j�{���pv����߮�q�c�^0ܸ���/r���s'c�r� ��e��tC��-��=��8h�o�CMJ_ͧ�����V��D!}4�}��q��z�Kɥ��6�bD<�a�$�>�O3Mf�5�n��?*���S�brCU��:��w'�+o�����-���A����Rσ��x�χL����)��XB��I`��%��I�W;�Y���9��5�AT�G+�Q����y,���*b�b��>����070�����'._�v��Zǖ����Ңb�(�a��YfNP���#��O>�N(@�2ֿ��b��ReCm����Ի���	\l�����������z��
<8��i�� ,e�����x�1J�%���j��gkͯ}*���� ��D<��w�p�L�	�J�PL��x/>Mr����"�o���pO�y:��/�BZ�c�4�	��翀OL�K�c��*9�T�����$]7mUB�F�d�Y;09��r�=zͻ^��gaaFƟ�kw�� a��e�إTG�U<&�x��+ô����3v�P�_���i�ek�;+Y��� ����|��W��-x�n�*-�EA��P��HN �-�˛����n��Kݡ�]�?g���C�dO����мe����ք���f�0����K�����9z�FV>���hJ�|�~�ab�/�䃸������T����*�v}��o ��`" �߿�U��JN�0y�3�O|�#�S� �iu�׳N�mm�	��ꆁ�9n�Q~��^���m��A#
[qB� >�6+��ੇmh[^U��T�C��
����v9���7>@�2�='F���2��Qi�L��:�RY��R�FZ@�������;ǩL�T�v��I~�}߃?ؖ3���$�QH-+��*:�� Fvp��Tr~�%s#�?bІ���lV��ϳ�<E#�yk	z_�.W3��cc�:��#��.�����L�s��0�<ٳ�#0�j@��w��>ެRo��7%�ta=k��iӌ����Z��h�a�X���"�e�ɀ1k'?�ݧ��P����(�1�|�)�Ȋ�����IZ���gL��R�k@�Qγ����t#�N:�7�Hiw^d�)u����S����2#u�I���9t�4Ev��������sQ8K`N�u��t��ԭ`8��Q�X��{��t�so^%m�-I;�N�j7ƪ��ҙ?jZd	UW��	�R	F�A�>�JZŨ1���&EH�Fι��Z38%z�n�Q3�{�͇
��En��t��Z�}�Yܹ���0�!U��/�3��y�V�'&ld�>��	k�ݘM���g�~Ȋ�B<=�T'k�y0���^������(�S~6�h�Nj����hQ'sQtJI,*�%&)������XU_�d��v��	#�$�_М͇�X�fY�&j���s�(QB)��T���q�%�"|,��Nx3��G�,T�̔^�����2���Y �1��s9��8��vC*;�ܽz9
��t#ۖ�{R7}P� "�:�.A�dei��pV�a�]B�7β��6��ŷ���w�Z?)ZZ�^ʊ�l���O"��5+z._2����/e�9�_H��2�-�5�L;:D��I��oZ���s��| �6*�è��X ޡ��-�4wW�A����{T@-ŏK^��.�� �k�^�h�,*V����y�9���;��Wn��ʑ�-�+lE,����/c'a/�^�a2�*��RHJZ�5�*�1���H��F�a������*������L����_��i�ڶe5�K���v��Ч94��/;�f�6���N�Jb���_�����R�9$����f�:��3T�(Xq
"�1x�?0��W��[�������(�p�4����o�5]s���M��� ��?:����9|:j�c������R=�a��\2����(��͞�Dџ_u'1���L�W�z�����#/Ɓ��#���D�g���v�R����ݣ_� ���R07&��������|
#k�W���ȣ
�骲�-5V���J �~�C�6"�t$QG�����+��:�c�Ë28�v�!B��D1z�X;q7�i�0���2O�����y�Xb�n{��_��:���f`�gU�[�)��粕�c�kGuw����-��Ղ��FZ��:-��l��-z���pz�Lr#&�~�'<��� qE�8�h!��S�a�-�%e���-r�v��9MH:����!��+l��~-�Z��şK� ����;@�;����]9<�U���;����c.���:Z��ss���0&���"�!$~1B�I���L#ӝ�A�n��g����+��9�����sB�]���]�Ԩ�?	k�G�Zk��Țl���4&�}��i{�B�P��<-<�%~�������E��������u��H>�p(��N�&seq��.W�Ļ�^���������ǖ,'(�?�p�/�;�Vf\�J#�Ղ�����#��<v�#;>�Y�WG3G(�ƻ!ׄ�d��R�narc�-��M̘�t�:#qP]�ZI3:z�z���*��m�µ:s��)�V� �*���>F3SbtӮ���x޸����F�%��ї�U�x��ٿ�D�?�� �ˆٮh�bBK@��y�U�j������ُ����ǥ	k��-Y;��h�U�_���$t���v�&)�h�����g�ó�=��2	��a�>~%�A���.�E�qW�ڣ%�d���Brf�#�(<�Ŧ]Wz��d��i�P3�!�ǝq��$�D�0)%~�X�O�a��w�m���z�-�M����lی��(�Sv�'fbK�DE��6��q.������B�lj��E��|K�5��r� �b��&Y�@�@�k!����5�\|�E٥�M_�'*��&W�<c�H�-8�%��'�D�5��n�h%�PED��F���i,�ܵЁ`����#T�p��/���� ,W�������K���o:��-fY��j��-#n�#��gF��S�.�Ea�M�1�52�t/�Z՜L	�����g�i����A���.�r]C�+5���߅���?�Wu���]�\�@�4_��="�؋��Cs�2^�M�
�?��S��e^�Z���C���R���$_�5 ��:��M��1KV����/a�����b@���@�)|4�����Қ`���`:�C�O���;z��)w�r^�b��b�ս����&���jڌ1l�.�L����{{]Wlù*���=\�3Z����bWŏL9���@��
�`ݓxԟ��+�SrKS�Daͮ�EW�[����>�$�����x�d���e>0�L�B���2ƴ|����z/���nZ�|�Ш�x�r鎜�P|���7w���Z�FAt�>�N�f�ǿ�{�k_g��]�]�%zw�%���M��o$�/@�E�Z��y]5	u�>�g�;0�Vq��ӣq�����٥}3Z.q!2i�z{���F69��8��"��q���R�]u�u��z<��0�f�!}Z?���HO��\S��������%�\]�B�\��t��4�$8�ۣ��[��r<̿wF��,wLF��`�'���ݟӤE�%�$�>-����%%C�;q1��\���Oe!�K3]Y�+�i��,�x�<��S7��gg�c���JjCҮls�_��x&�k��bp�WX�9z؏}n����7A0'�R[
y���.��Z�m�a̩�q�g�j�Z���IQyMw6r���C���oC����mw�\��g���֛��w�Kf�;�ޮ��8cL�ُ2*Ӳ1n�٠��4��8��`.ݨ��~��ǂ�ż�Omֳ*ht�4��`.����bK����Et��ř��#K8@˜�ô�,U��!�qK%̆����@f����m'*����V�H~�%�U�d���4%^׮$�]�yu�9��dR��%?YH_2�oA�#����/qaƬ/��)N�9R�B�3�u�j&&����b-�<�W���/*�>R���M4#M��{��K���-��V`�;��q�wX|�[���D�|~�C��Jh*U\�p ����ِ���nQࢧ������	�]��73�Z��i��*k�8xF����y�4auS��d��'����+����'�x�;� ��WSJ+��)n^�?�5T۬ �ѦN����y����\l�m���8���X_��c�P�I����%@Ŝ�hW���>6�pɿo���z���9RK9X��|��Z����\�����^®�ńSy��eb�뙊{�K����4�_M!f x�6n����'a��dױ7�Y�0tnh��|�\	9��2�a���0Wc���y����EHY�5�+�-�}�&�c��ʎ^HoL��h��L�w�àu�4�a�]P���\ܾ��~0�3,B�N�:�l6�<ƅ8w�4��.z'�)�'�s0�g���p��}��?�hg�����q��r��a\D��=��)��c����[�Ȏ`��H7��#���!��x.$�]Ȃ�6�R�x���A+� Y��9��$M�ˆ&Ȟ����E��۵kB�}�7Ol0[oO!
��%Fznd{c@�}~�:��Cȯ�L�7C�	U	��jQzd���T�]_�t�e"�?c��\�"��Ȫ[R"χ3(�zu��CEx,^t��ɅoMȭ1�t�s��8���J6vM�#S�������l�,͍�K!./ �H1��)]��:;��s����d8��V���7@MPz�V��qn&VSؔ��	w���� ��H?�i�0�@��#���&4����BT(Mk+��mҭh_uc/ZT��ە=La�����z�����
M�����n?�p
�[(��ĝe�q|��
;��QoTs����oA�Q*2��$���f3��k����� &����균�p_�Ud��d��N5午�?K��ݨ_l�Ul�a�TqM�
��B��D;�x�;�.�\"v��0C�k�u���uC���u�ۆ��g���H7���!�r��x_ ]�:dZ�#� ��@غh#��Tn�����=
�I�WhUV���[�����A�e��KS�,ī.��!�kz鯥[9��Fi��3hD�?]�mF�{��o��[x���ͺ\��p��v��ͨ�3���Ȣy�%I�W�)�)"y�/�"V��+���'`� @���v/�|��3S�|���I��*8����io����l��;h�3���nB�أ�R�е1e�MS���m�VwZ]R@�^mba�Z`^��y������XhZ��4n_��C�����[u!��AN�hw<*���4*���g��)q>� O��.<<	�I%l��F�{W�5�$�ֆ��
��XA�%���~L����B�@yG��o4�a�B�4�?���e���#���Onx���`�$�9t�KЬS�`^�� ����BΜ}�S�f<��fi��a�>��ۇm���ya�JtvsZ�4f*3��l��%pЫ蠬-�m;�@qT���>,_�XuP-�p����(�UPdV��]�a�w��4S���{W���;ZX^�� �NҍE��ȷ�\,4^�,F�s:Q��w �����jv�9� 6��J�lB�-3�W���b�m:�2�$VΞ�����Px�\�D���<)��Ƌ#bC�:�9�I��@�+��|9��5���S�jP�8�>��9�ؾk����D{A0%N���>��#iߎe�^."4n�m�^��@U�@�8%���"��u��o�u-[���	'�BԫQ��Ḩa�¿N��y�H�^����=m����5�d��r����L�����?T�S����_�v����+yqx��*�P9O7�]�_O|rW����W �HS.�^VK�U�����]��b�%Wy�Ȅ��j5?��,���֪]͹�V���s]e�]IV; �J��̭��ȮJ�s����/�*mm���Z5���H����m��Y�rv�dڎ��lk�x��^�u"��\���U0[2� \�O��F�qx��6�vݕ'OV�A�I�Fa�EԒZ�����)'������6�U�q�2�I�'�R,��R�[�oz���p���=`��*`�e|"���א��S �e��;������x�cm���c�3���2�t��x�(]JH��g��ˇ�2=�o*|H���&�_��B�9\>�D�<�gY��B���&0�Q����~e��
"��%F��0��K���~z���A��t�����R�O��/r�D���tO$�OfxS|Q3�«�<��+�i;�i:wFa�X<�"V�&Ȳ�p#ǁ*4怠lB/VP������i�R�����͇�}�mЦ�Ų-Y[7gN�6�㫿�צ�Օ;sWLd�#=���KhcR4yB�AjDW��>�B.���!i󫓢�}�����'��)]����V���ɖ2,���:
�.g�oCɫ�ҧ3�ɥ+x���<��b����=��.I����(/��ʌ�5�r������;���=½��!h .��a�Z��|�`*�[���J�Ǽߘ�*�h��f '� F��t>�@<�ٝ������2
D/���u��+O
�'�1�A�̧�me͜ߒj��w�2I�R��Y��=�x3*���̧�y;��ӫ�
1��
�}/d��}�F����`����O<�6`_�A�oK@�E,g"4�����2W�)������\��i\�ÏfG�vj��r����;�D@�l� #����{3��=X��Ԃ�:,��w�rlX孛( 9�NB��#�ğ�Nb_��)�'�E����FaK�,�>W�f�� H��ﵩʮt�|����F�(|���
��M[�ѳq)FaU͉�{} H2��&����9��-3-���$�<x�ahk�c�� ��WY]���o+��Z6	�D�b�
�bUi4����H5f��_1��]e&�7�㕙b��ОQ�������o�6.:d:�$m����Hv��E���Ư_��z8O:� �^��x��(n-,0:� �L�w����v=�ss:ۿ�)���&����FקPH�S�� ���C�?w��?+�����;s�~qi֬�x�L��n*���29:���ƶ�\q�Fz��1��UǊ4g��M�as;�s����?8�H&����򫬋���V���h�R���A_*HI�B��S?p���v�[�:T< ���17�m#ɜB1�2L�`ʦA��F)M�3O��NoG�؈k=n�+NF��J��Ig^������eԁR�	��LZ���G�sL���_�w�=��e%q�f�M��(��4�`��CK"w@I7o���d7���}J�TR�����*25䬟�T? �]/����p�C���׏c'ί���~#�%3Ե��,-fڍcʳ��h��ѭ��I�-�x�ZX�i��������<`��P���E���ujP3;����%太�6�4���r�V���(�2�z��}��گM7��h`�u���~��
�ǥ�e�����_`��O�N3�`�Jg�zہ7�,��[��=w�� B�7�t7$(j�GRN&�w0s�Rq������q��__��F��k�W�O-#�A5�`����=)C��5�	�wJ�/�B2 j_�]rS̀����#==����'�@�����B�ovB�C�KҩB��2����������k��.�"L����]WqX�Np,`���G%�F\���=�o �RS�O�ZB�]�6i���е�E��+����x��b(� �*ŋ+0���*
�X���f����k�pQ�}�Ӕ���[����t��fld#]�!g� �0� ̗zң�7�����dU�j$���<�V�~�����5��w߽��F�]��HنтLl�1�ұڿ����vh+�տΔ\����j�Q�g+ǡ�@��<��ٍ�߭R,�,a�� Y9�`Ú��{��u��#n̡�_���#�V�:Ͻ<?���7��V~��)�]n�����"�����?�cd���j���t�
�ZXT��Q�J���>�<�m	�nd�z���ۖ�bnШ�
�R�Q���Ձn������2iN
��V*z������@��#Or��G��L'���B�H����}բ��x��������mE�Еo5 X>6,���2
{���E0$Z�W��H1�7�j7��'XL��!}��O6۹�!A�?G���m�RL��P�vx�mF����V��+���\L�M�1_�a�)�v�����]�p���O��^W;���<O8f�V�V	T�o
E!��@����ۨs;�r�tD\��T�@��]aD�� ���+��/�4os��J5�n�i���Ix�S%$	zF-R`;1�-	�8Q7�.9�a�c�D��q�`T�+H@,vH�
>���$��RV��(f��-�&AHJ/�.K=�����tgu�1�8_B:��M>vx�T<N��|W`3��6��IȘ��j��w��R��G�������+�?oD@�+�	^���O��k��������*2����"��ߒ<\9����؇Q�S��]�"����H$~$c
�:��~!�-VĨ�K���1��*��E=P��G뵥+��aKAT�q�$�-�ȫZ'`4�\��e?�8̀#E�{Z�\�u�Aa��&�wW��S-�&C����ٱ�!ٕV�XR3��T�|�� ����*X�xQ���
*?/��vA�Ն��fX��i �n�J�⑂�o�K��1�1󁇆iZ�^?��ꚜ�>u�e��R�^Q\�L��u4�ه[�M�����@r-�K�;F�;�[���O���a�3;S����2_E�O_<�t���<�8׻�E�M\2Ŗ�6|iz{;�U긣�q�5`�>��<��H�iZ��w5�yr��in�Z2�1.���C�mԦX6��0L˄�ಊ�Ee6��S�M����O��H���͸��J���Sl�+��e�����m�A��=~�W�2�#�U�7H>3�������F��k%�	��\�lX��w��>b�?&�<f�Fn�!p�&w�'�����dt4�)]y���U�%8�L�7	gV���R7
P�{O��"Yq��3�i�B1�3�(΂:Ǆi/�������Mk<�i���jԩ"y�"��I�U"u��z�+�Ju�+T�τ8��ܦ/.�%b|yv�`��	�
���	�zGU��Z����
I���V�:l�:h� ����T��l��ʅ��X��E�i��x^�A���;;{Ě�%��W�'�F�{n> �n������:�1��p�=*$��G��D�N����O/��BC�Ee�!DX�i��5�M�I�����M��ߙ�_��.�X#4;��+�:���BH������E�9VMi�����
�D�շ����њ$����ۅ��N�M����y�����%Pb�eF�X�p��mJw�^�v�!2�
S���?Mv������wZM�Okȸ�n&z8P=t.��ߟ@��mPI�ڽCa��LgI��&w0E�/QuR�]��CC��� ⥪�.��}X����Q�Y��t�Q���UPř�vm�h�k!�[	��A�Aft�h��Յj��cm�D��n9��
9�����(�P��@A���dss�����F�F�򟰉��C���A(Ěf�Y|�M<PtӾ���|��� m���/��������/Ь��-YΎP����k�ׂ$B��%s�X3��Q��ݲ��sKDZH�-*��}��.��us�7��b��9��4�h�o#��Q�>r�</����4M�:��9Դ���� B1�{#32
7ɖ0�����f��JF��M}�;��/�������.J�lQI9�W82Z�����̰���EOg Rf��$	.j�/�P%&�ɵ��������P�����NI�dk�\O6 �BZo��勃g�o]�4��XbJ�H%���x����g�"bs�:�Wl����?*tpDz�۹#��{��tfk ��vƌ�L�L����Q{2-��kQɛ���>�x�Y.�z=�>]y!���y���I��|cQ��=�ֱrʑ�1SO)Z+��3����C�+k�n���ʠ'��ذ
a�~E��4�����S�i�N�=6q��|3([�N��s�jF�H>�=�!�J\DըP I�˫�U�'^\�^ u���I-j������L@*őE���ڂ�^�V�d������S�f�9�ᕘba���dLw�����3|ù��K��T�@����qҾ���[��q��D��0`WJ<���KA���=�+	g����,��Ah���6�/|���b�k��U�U���Л<B�~�gv��5���^O�}��O�H�c�v59[��P��o��π���Q�(<}Xs&���
c���L���ڣN�