��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���NL����ʇd�2e����� G��ME|f�l�(U�A�<4�m4���u�*��n��_�)>�z��?P7��E�%'��Q4�su����p�|uLr����=��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�O�5t�"!�� �RY0�J���$��x�+�D9���m�P;\�<�"g�W�	x�k)*���uj~��H�wLj� m��I���%�k=}胄��<�v��J�޼1cS�h�~��X�?��PR%rs��8P�W��F ���-�R!��鷧+�7J��j�f�ͣ�H���5IT�������B��+���p�"W��j����4t����O[��:.u)�-�)�u~o�~\�y��Dbm[CN�愴Zל��<�S�Z%�^��^�� m(M*��'u �Bf�[�Ԟ��"��w�0a�Mt��#��zu�<,6��-#(@h����s�;�F.��1ӊ-�����qo�`���lˊ����+$�-�"*.G2�_�=�\�I,�)����RG�����ܘ��/���Z8
żJ�K5��=I�	B$�X�w;!C���a�E9(��n�hY-P�UȔ&j'x͡4�cK�� ��[ҟn���Xb�����W?�F?�E	��|�5��� c{���5^Ƴ"��~ �j���ؾG81�8�?t�P^����nW�r�'o�kP�;dt-��R�D��G@t7�x`�^�LTCt�m���8A����&���!p:x�u*��X �:�H0����o�~��d��N�p���*�_<a�:t�^
q0�t���38PV�#��,�p ��{�	HdeH-��e*�h��XYCa�]P��z���t.L�s�	���&������
���G�%KE���k�1�,龟@�Gx�sb(��ǥ4�����'�Z���}�6���s(�Hg��H�*���#*�(̚U�}�h����ZMX���WU���a=��Q!<XHҀD����J!@�*eS©�ۛ�~@�zm�FV/yS'y�ՂQxrI/�\V��T3��{C�X��n9��ّ��P[����&T%'&x��
O��y�[�}^>�Ζ���t,u��!X�~u�̀E�6��xe?<S��Ɛ���[,p�.��F~l�ެy�&�|�hgNshGh�n��+�R��� ���&���7�@�le�=���a�i=y��?t�`uE��e�^{��V�.���O�?V�6���D�r��a�H���,�Sn�Y�߼�I�A�ū�������`$�ܯ���x;�Q��u�s�
���;Q�C���9�.z ���u�l����D��#���R-�zid;8^<�Ja�r�Cٌ%Gw]Έg�2��ߘ�T: �:���Jk�� 0�!̌�cmo�(�U]4�P"cu��#HU��'��w?����b��;~m-��&��D�b�K1�ce��?Ly�.��͐�5�7�	7�a�ˣW�s�^є;9���
s���fh��	]�=��X�\�N��Pi�i���ş1zⴀu�-���㲧JPe�=�Z.cd�sfm�[�0
-El��E,�梣�/.�PnY��`X֘�7B����R�H�?�{m��KK�e�s�*��[A��ȵ:�+'��7�����;�P��h�FBC>W�5���X����6b��K�WΣt��0+p8�3���z��e��zA����a[��ɴOq/�˛<l�t��h�ue'аf��j�V*-I���g���,5n�8p��p�%�����I�N�3�Bc�$C��t�*h�IV~P˵�Lo�C-�NZ�	�	Q:[��l�U�aѨ�	vҺ��=?E͹�Ew�v�:0�����6��a�hp]��E��V�"���i�K&��I��OT�~��4�)C���n\U�����n��	��?��d��P�r(2�	|G2{^k��e�f��}���9�����{7��Q�@t�p"�Ϊɼ��I�M@Y�4�4	���p�����;����Ml��*�Nר�j%rq󂾆��2sA�h��Xʯ$�"�k��B��S������y����@���Z�E&%�/�����))��!��w��k�H�����^s�O�,_��}���ҳ���ћ!�##�n�����s� ��x=��:>�
ю�����_6l��E�Yo�����`�_y˴��U\S�R�c�]��J��v��萶�YlϢq���= p�3��Ŋ4���Z��T`�*l1� (Z��|7�ڎ��:&*!�O��w��c. Gv�y�bX�g�������UX��o�*�1�_�B�영&��^OP��q9.\��$J��`)S�$�c��������\���#ǉ��C;�(��ĵn��6Q<����Ey���VΫTS��#�0䳬B(g�CH�U��<k�ːԜ���������.��D���$\PXw}���-�嗾,�ȴ��%	��z�J�]���oN�
�}��<VH��4�{��h#����H��{��?]L9�LT�H:�?/��!"
��v<����ّ7;�~�R5����ҬN	b�	�è!����5��qߔ��ц��r�����v=x���FY@v�%���6�d�<=yH3@C5_� L�2ѹ/�7*/'�t���&8���V�;�NC�o. ���j�a� �ȁ1[�k����:OH�TF=��|k���.nC'(R��f|�KX�#�)<B':P0��i_i�ox�hHn~�"���!o�q�Z����a�cб�H�bI S��D��8}�i����3�, �m�EH��� ��,�������uRl|�h����ԇ4>)�Z����T��M+���MNkK��5�~�'�Oߒ��w��;04�!�k�W3�R��i`MdAߴ�C��˞q�Y,����{�Y�<���xM���t�D[8����!���+Ս;NWG9@����?¡)!|�D��0�Kڄ`l��1N��.�0�S��;����DX�����;݆�P���vK��FQt�R� v�>��r�j������#�|�
�rO�$!��>��4	�؈�� �1&x9��>#fݨa0����]���\�w�omy��BZ�����U�ӏ��Z3�b��ߏXV~�� Fn��[(�`��V��X�sXo�l���=�*������8���`�w�P�9�Ff�*�����YY�l�E��3�p:�9�U���h��������F�r[��,��/DpQ��_Nĳ�fJ>�P��o!r��[p�:��B���Q���O��rD�Z|�O]���79����H���!��^�?S3B���:�����iLCx<����|��0w��M?�{��h�U'��`�x0��OY�~+X���<����e���eo�O	N~�(�JpȽȬP��s3��A�6�i��jƿP��ƌ�Y��{^3Z����cv�0�4s�v�����$zFI3>���0���a���}K�R���$�Q�=�S�K=��c,t�r��NJ��.k%)9�I���yq
ћI�������^��4�C]��8�Cd��r�<��)4?�~��zwq�E�C�'Nw�b�#�`�E�g0q���B*p����/ۧ
V���|�H	
Oi��8hCҢ�Y��R;.����t���O��Q��G��|�w�o�mp<���f��ba]|���S5�P^|�IM7/8
`�/����Z��Hᯗ5WO�@ N�d	�fv�W�yZ���n�nZ��x��E�Ķ?��] �6,���e�j�e������-iICm��������4�F�|�z�~N8�a0�T�f�r�S7�Ժ��W�^�(̽/����Mְt����لGkVP�*�{��7�7����L8f��Aג>�ސ�lB��q_%�pP��Y=�ċ�2���e��"� ����t�	
ǟ�/Wf�Z���;Q|e�F'���lM�T0��-��$��I�Ӆ��������nj��7{�NZ����x�i�����".�����"0��R��&��}�s����O����-"B�3;¾�,n��:b֣X&��1�������F��)S�
������	3�`0��
.��	F��8z��Q���Bv'#��ɲ�8�p�٤\�,\U��H
��b\� E�h��>��*�a�������dNW�=��F�O:!�SMF��ǝ���&�/��(�P9��ѐ�/GPO��ȃ�g�MRƖ &�z���ɐ�4I,'m ���N	E�MJa�����W��j)����M�<�vqe>¿f��^g�{��-ӝً^��![G,�4 3�)���Adτ��Y]?�t��f;���s���->_�d瘋m}�|���|-A�+�Rn)4��`�����{�.��:F.�����_�� ְ��'���q����v8�� �$���j4��^�k	�Ƽlm˃�N_��w����蒸�uf�~L�qxL ���7O5�?���wb	pRw3��=�j�~*_������L��P7���9	����Y\����W��}��PM��sEOw�^��|�]���z��� ���M8Y3��j�m�r���5J�b�4jA�$�d�t/wN�ЍA.E���*��鑩n���!g~�+��x�PЊs'j^����44'Q)�ƜڰgW���S�ۗ��*i���@\�IH�h��/��E^똰���3&�;����8��k;����O	/�g�5�N)+'�סeO��-��ƪfYU'�~���	E��L�КڔV�_�~k�������3���ןsR�9�Q ڠ:P"(��v�C6"���>��R��#�G�=���6�1�eJ��ڲnj!�m#YP|\l�Rݵ����I��woŧ�<Y��6?�6�+w����4 ժPyu�I`�'��f��=��(���5�jL����c��u{j���V�X�`�l�Q\Fc|���W@f�<ʋm0�_�n6��0���t��[��v2�C�n���]0�v�@	�2� տDA��X�������*)�sI�[Q �!6r�Ӳ_�o#�ғ������[a�eN&�n��YG�s����h�JD�p�S+�?���:��8h0_�rs.�܃�����~��볥��w*�!	$Js��* �T�˱�����w�HTr�錦f����ӵ��ٚ�Q(���������n`�,m,��[N�߹Cl�!%O���=	fy��P&���,k��G��ŧ�.����́�ha0�^�oa�S��9�t� ��6���]�N�������Ԩ=�b��|O=�g�g��+��t~������H�/$�S;'���6�..�(O��}�����⣰<	*�|��E�e�������c+�:+��A'{c�O�G�>�н׵w�a�ta��,��9&Mw2�C?��^���k�f0&����ToR��y|^Dx}�2���h�]�@������ʹ␅����(-,؈��G��: ����/��ܴ'�Ց%	����`]�/�D����p�|�aqƶx��б�G�U ۤPT�E�Vg&pl�\���2�������>����H��O�f��\3����N.})�vêvy�< �Ȁ���טU�U�4i����2^��M/ �I#�||�����h� ��ڵ�����h�w����O�a�~��80��������E=���,RS#�(D���<��(p�R�>��)�]Ϲ��*����?�)
ǆ@�
���l{M�K���+wW�,�/sYm<�����clsL�.�w�u~$�p����.��?^+<�Z�s�t�S���(�?��-�i����1 $��(c��߄��v��D�(���-k����'�/��6��\/�g{1��g�mt����:'��0kW���sR_ ����s�xm���@`��ҫ��L��mZ��g�--��a������ڦ��T_%D
�X�P=S���"��%���'�k}��cj&[���ѕ����RЮ�9��F\�~�Ԍ�Y;k� h��XB���16��Pۮ��d�ۙ/�k�C-�Ǹ�Eԓ`UE��G颠̻��˳�3r�[���!Ϫ��Q�u�q��?z�c���S�t�2�O~�ANY�k}�(*c�r���$)�TjPk���k{�	X��ν�30�� &�����
�|�_AaL{X�wZ��YH	
ǅ74LHbF�����l���	,�A�Ԇc(^ڧ�J���gx�Y� $z�T�;�=!J���y��� �_����Rc���4��G�F���)�8^1�כ><�l��k�g �ҡ�B6�k�r��`D������y�3�9�98�D�K떇��;
�lɽ�sF��=$rJ��q���VP�)O����5���%������+������#��L`��,8��Y ��H +�]e���j��_���;��T���Lݫ��
b^ 	n ��s��E@~4S6KtX�Jo�"r���C�VQ�`�'�d��Z<�l&�dc���˭o�,�\ckٸ��{9����"Z�xHo��Y�*h]뵝ɠ�=o^��y��@�70;�	�P�$���]K&��ָIL�8��ҋ�̌��Л�i�Ay�3��w���Pb�|#��zW�_�6�"׻FN�P�M��Q�{��c���H�V�Q]��i۱��[`� d�6|�rw���u�ș�Ƿw`Yr�\E�ݒ��D	+�3���,�շ��Ki�%?����4�ZD���؍�z(�c����WC^QLQc�,Q��bcd;�tI�`h۫`J>,7u&��WF��}�M���(�=T��	���t�,�y�
z�t��/��WAڲ����]��E��y�:Z���?����d/H�7|��t7M���fg�:���s:H��7�y�;��g�����:u��,�|���'�!���!����/�������`�m�0�L�n�g�S	V�r�K�S�����6��]c���\��qǢ�f����t&IHP��3��de����@j� ��b��k�R���ؿS4�U7�(���[ͅ�@��7R����w��.���O��`���l�8h��U�8#�BѼUQf&rcP�S�=Ge���|H�+~�n{wE:z蓢Y-�
��tA��M�³j������o	Ba�|]����⮢.E{;o�Խ�F�D��5�{�4#��]���7�i��M��3*o�L���2���ō�WD��I��{w%b�",�(�n�[e����}%��yhnj|Yۼ��=�:ۥa���4��u_%�tJ0g�"B��(�{Oи�� ��L�S�8:q;��gv��Ѷ�FHx�N�4k��N����ە���91=EM��$<nZs�
x$N>��e���q*�h�tly��=�!yȑ����J����I����k��.!�[�L����ΐR�s����!Z�b���4A����6.�o֝�ڌ�*۴yk�*߼hA{��ƌ7Z��G1�V�fV��.AU��n����J!PӦ�k�In�
�U���e"Y4�i�yBn�TE��U����>\��&Kv�n�PP���4$��y�k'DtV񸛨5f�3����2reyk��UK�1u:L�0��P�bb�Iؓ�/vE.���C#b����Gʞ޶���Ĕ��H���@�&��6
�n0�����!�9=���J��)���\���vW���?``K
������[�&���v��ܘ�@���E�3j��g�*��x;z5�ژ�����Ɖ�Uȫh���x�>����ְg����s�4Z��bH�2������-J�S��2u��m�'iG��>�Re���V�'M�� AZ��溋��-�z�ޖ�3g�����5r�}�g�<kLΎ����q}����X�Ə�ӅQ!/�\a�]۸M�De�r�El%� ��)Ə����Иa�>�Jq�r�|m+�p@��v+��C�e�z;�h}���TPŹ;��-q��_�ǈwp~Í�B�/2�����P��h�&��~����\�0�����ݨ�	H��J͌yPG�es�˹fù�ϸ�LW�A�lO�r"K�LJ����L�'1
��Ϭ�Y�%����>p��������L޹��g�GH�頷��n!u��Pd��H�ﲅ.���#��t�\:-8��RgH`�R�$�g�]�C�cP��?����K�.J�Fw��O�V㚭�R
�;���m��J�x���V?Vq��t{j���_���}n�Q1t���
��@&����j��H�����lT���"�;=ˁ��1�<� i�SX�q�ƕ�Lu�f�0���[%:,w�����	Y�^շ�Q�H��x���/�#��#�4�u>�T�)��(��HY�P*B�Ӂ��tF.�S�$h���~d�����d-����֟����mU	�$��F�V���Z�L��6Ư'����I/���(lK���|CEv4�iLOY�������uQ�E!b��ظ)�M8���ש�r�܍��w0F�F�[���)RY��=�87B�����s�YplE�uǅU���d^�9�ַZ�1�&a`!�3�_×��x�yOz��	�)O�0�����H�=8�+��O���Xw'�y�r��-l'[�X�w��8whJ��az�D�Mh4/�`�k�_�y��y��*����6���� r����2(d��;����F���O����5�
~y�5C挻�X
�Nc���Nj�<��WV������4͟y�E ��>�FL��gU��b�Oq��O�8�԰�\<)��{�o,����ME����p�U+1f�G}�h�]�m�]9�|�L�,j�J%�&��=�+�-��̦ 9���Bl�4��*(e��]e`Q$�%���Fsg�!i�VQ�q�Z-zذhK��ژ�L:�Gi�����s���Q�I&l�כ�W��kK7T�n���dlb���¾� ��Qn}^�<@[�L�cq���#2���(*��(}�;�'��/h-�6������8�����.����+c/\��]|β3��q��p�(Y��lʝ��E���g�:g�@~p��.br�5-��O��.B,7��P��a���ц�X7!Ф[,�h�Χ�7`��	�xJ�</�E�&Hs�oJjDb����,�h�a��2��.&(�6���M��ׄS���,F�xr��̏0g�k���N>^��  b�Z8��I�:P�6�������P�i05�?cOx�����B
�1�\��,�ѪP]�Bf��\3=�#C���~hG�W�p�3����\p�QU��D�<��Žu��Q�-}�U����;ol�%���UZĆ%c��S�.W�W�
f@^b�S���N�T��͵�=!=�E�y�[N|�09�Uc�E�|a`�x{�� �u>���H.e�.�����apq����[ҥK��f[�� NU�~�\����.���]���,�r�/`��Or&nS��iá]�r����m?���% �[�T̙����QvPV�Y0���9#����-A9�18]ţ��h������L��W]Թjk���q�^_�C���Ñ7#�<ݪun�8�V�Hu�(`3���O)9U?���`%�g�x@O�j��E��"���{�4�g&��DE��k�*Q6W�iRs���6y��c��$��K&n��c�OsK�9D3~�G?EV}��Wآ����M��Nq0�A�����[sDV����:��1(����%f;���I�F���#Aܠ�zM�"��z��|��1��a�D�;=��2#�^�Q@i>8lv�Y(O�`��^��uM�����dw�!(qE������$�e�_��)"[3{��`$�"�� l6=I�Z�o?-NgI��Ar
4nB��f�������b~]q��֠�j�<�،�b���V*�$���S�G�X���VW��̀�1"�eS��,�𲥺&�2�?���p���@����o��E�vqq1E$h�S�}�ei����K���8�{����,c�Q�:��Z�y��`M���{�P�h
�#�pt~~�`K�z[�c������k�|�
���x= ���LF=~^a�n����H���FK��� ���qL�[��MF\P׍�� �|���h�DA�_3��pT@U�Xd�!#�Z)�`L�3��Ke,��v9Қ
ļ�ߔ	��X+�	�Qc7����?��M�1ȃdw@ z��޼�T,�n��Q�<� �ẅ�L�FV�~�4�W�!w�s~�){���%LL��0�f��J7��Q����8 Z��
�o���?Y� R�Y�ܭ�@�z�W�U<�Bo{n \��@O_�_e>'mfC��E���3��D3�S���p��Y�s\��,pJ�2�?�ٸQ��_^��l��U�_ESk���J�~����P�N�O����|����S
}=�4r_"�����W(�������Cdun�3��}�~[�͗��-` ��cL�a�A�mjZ�$l��Cc���6i	�l�=!�8:��`\g�s<�I�����{9�B��ȃ�����(�A��:1o"�L}j��y9�������l�߮:$�$��E�0�+8�����,z[ig'�� ʔ6Ř���W�Ad�o?t�!@�)��b�������*-���i���R|�[�qpQ�6QI&���s�n]�i�[�τ�TuD�A�F��o��P.	���B#a4�$�XvLv�6���w�>h����BD�Yt�iǥ�m�i��l-8p���2z���T�۾��=��\ب���W���/}�E��^��4�3��#�ve3 ��%����0y�R�X ��b�[ ��))�)�#�_*�OJ����:Nv������,;��>�.Uԣi�QAD��6��=�d��g��2k��oV���� �^J��ʃ��2F|+Tm��5��ڞ
��D�H[�oQ,�m'y�^�nb�M�Z/Cbи����� �1�m�%�\u%U�_-����e�6��S?r6�0���y���4iƼ����x���ZM�}��lY=w'��ź�ۊ����t�%0�GĻR��S�L4�{p���&<�ދ&�������������Mm��_�.m�Cȇ�R|���AJ)˝]l��ri1`%�$��
NL?Y�c6�6e[�8$K��IF�N��L���������*���8G�	O�A�n�Qz��ef�t0�йs�#�ÀVѦ���{�Y�긚J���ah���p�q����&D�0SL�1��Ӊi�K� @hXBv#��o����	$���bٟ
%Ob�|3z�`C��0� �@�{��q���e;��@��Q< ����Q�C��e�/x�@�OgI�J?�DT�Eav]:AR/ݠd�ev�pMA���]U��h��~= J�P�0ma�5Y�t���&�A˩�s_�tS�,G|7�>�
�/��Zl�ه�5NP�$.ۈ���-���Nwe��E���P.�#���^Lr%N~ ��X�Y���G���I)����t�s4Յ��ߢ�'y�S ��G�7��W߱zr���' ��k��F��O���s�E�kH���*mظ���lᷤw����)������� �u=����V�P��i��O�2��z8޼Rf�EN҈�sΦ�.t ��vWV�E��ڮ��̒�Y#kD����ii���%!Ce��D�A���ӻ���j4V��֜#��j�E��Ȣ����<����۶|��^)V�0ȵ*�CL�׫����������us(\Au񡹐\�H!2ѣz��e���y�4�aw���fSVM˂����Y�1^��ƴ����iatX
Ȋ>�)܆�����A*K�q�S�Z�=3j,X/b��=�G	je�5z9G��F}|�x�#��o�DΩ�PdE�f�H��l���}N���>ßf%�d��/1�PçL�����M��O�zD)H�myE_EW�cY���[�|G���\��ifXy� G3Q���]�����[XO�]���:�BC�bg|h�N�²@u?F�>���`��v|�fBκ31�)�`�n)��!�1��K{�a��/\�È�D��IF�?B.�9��6�}!� ���	<7���kf@d��
r;bv�%���|�n:|g�Wx��&��;h6�£<}�Hh�'/@�Uu�!�PO���x���a\H�ж��p"�'}k��
�.��:n�7GGM$�:`�e���[V���Ծ\*��'oMly�
%ⱘ=�;-�k�5���LI x3���8�'1��i�o��s���Z�y�v~��8�����U@
���d)4{�|�yު�Y��i�1n懮!�5b'���;ag���r�䄰�jb{��G�gH¹�N�o�թ
3%��|	�!�P^�
�%H� �%�:�M\ֈ8M������k�������4ܟ�<������p�CWZ�uσ��i�am;7
����h�Be4�,��*a^�mS&�uJ���Q��Q������R�����ō'h���#�,���zb��ȯ\�$���|dT%44�����t��#��/����Y�~<9��Ti*s׃�zrƩ�<}�%0�����#~��)t���Ԛ�?���&Bs�-9����8=�9,IF������P��(f������?<�2��b)�A[������YP2��cFt���n1�{��lH��z�v�I73:_��-G�9�!���@�e���t�;�KQ�ó��q�9����	�E�27A2:���?�\AvḼTW!R�g8j���|]1�T��u��;^���&.7 �"91�۩���2*�|/n�U�۩ayf���O��E��$���RT���]0�3`�Y�iq����5���3��C�j�$X�^̹�C� dz�t��@GS+D��^�����`Dg[�5Y&��-��	5��˗ѐmM@H�E]˺�}p!��>�y�R@���Ӝ��g� ��*Q��pt�3�������c.5oA>����kz,#�?^��E2���qku�O���9�o�h�y������TA�1?�](�ľ5ɑjtA���^��$��V��XXuJ$w7�,F�:�0t�S<�=ުA]�H���w��OA�!zǶ�9�KL�����0�_fY;5Mi|�&l�oY��jY�V�AS�BmB�������w���� �>�{�f��9���gq�072�g��ҷgo7�3�d�L�aj�m5���yo3�xL�V�S���N)/=�K�M��Ջ�����?`��:W	u/=���&"�Ћ"_�ѐd |-/Tc���×�p:+/�*6���Q�溢��p�j/kyEU� !���<�D�v���z��uL��>�4�/�Uնd�k%s�[�L��-&L��!����әӣ?��@',�����S��6�[?}�S�w��@��GKvw%Y���D({h��Ԑ��J)Z�&��� �"�F����Q	�_�Qbz��� �r����.�8���"��Z�ْ�\��K�dׂ�ctI]�]��
il�?��*�R�\jz�@�7n��ld�-x�P�n||�-�փ�9�2��Q)�k�fϏ��M+o�I@^�����s
�"�@�č˚V�����}��A$F�5��wQ'�Ae�����W�o�����C���"l5F~�z��7PxɄ�Md�B۱���y�0Y�� ��J&�N�}�:�iK���(ù�^����bL1���<Y4�w�iL�M�<�;G
x�VR��|͖m��axL����A}��7�",? L���VN�JFt6���#�#�R<n>�P�b\F4c�Sj�=�e �R����Fi��b�4]��o�!)��8׭u��G�\eƅU|Y
YrOu�.٨����hC,1a���߳�9�n�+=6��I��t�Z�e�¡ ��I�~��;S��rg�����(�ڞ U�<5]��d��T�?�����}ܘ�<�Aqʙ49Kn����e��Ʀ�T����ʅg����ͮo$ ��/�(9�@ൌQ-%b��^>ݾ�y�9�7?fbF�2U�� /FxD��r�����N1,�2;��=���"m-^�r$�
#���_�s�	R�?CNu�*���B����������Si�uEXoςN�䪫G�(�;a���a�Ҽ����-@K_'VO�R͊'Vjg��$�e�%C���@0�� ��?Ă�?���
j�g�y�@�X�TF��k�c�1j�(_L(:�CPB�[`���g������Fh}_h�T-�[��4�Q�=�h�n�ob&�=]?tb���g�O?���r��d E��E����7W8~�f�U���ҍ��[? �iq�N
\�q
(F��l}G���&|�`a������h}0��BJ�N�?%f���K6j��;ڄ��%��7s�{�!�,b~7Zr�wþ���|
�}�;0�W����A��>�{�hx�7�N�8a�����A�l��c
&��#兒A������=d/5�����e"�o{ _2�Vfp{5��ۂ�)�:M�K'������T���>�ӝ��;I=l��%�����I�����o�/J[��ବ�!��Vf�����)��ڦ[SPԑ,9>����c~��8�gp	_��8,=�3��E{��N����B��V��tY��/E�62�[��Qу-#���%�Ig���/sn��٭i��E-޷QI
��~�v����9�@!�c��?�����Mj!�6���R^ߗ�D��h6xΩ���+��R��*�wA\��TK"��Hf�k�5�	Fu؂���g���Њ�2E����.�e�v�:ڃ��9o�2(�K6$a��J�~���:q�3��6˾4ň1!�:���/`Y�zVv!qYC��EQ���|$�o�~kA�e�ciO�����AH�K��y��i�xxs����ZR�54�>�����<�qޚ1���Bm���ѽ�/o�k�㏘��@X�Eu��MH���'}y�sm�Gvd�Ցi�]'eU
s�#�;��`AO�n|n�}֮-�^����qAX��J��#�R�14�їF9�ÑT(#6��C��g@*��֖ �'�b�4�ݭΠ+�ٕ&�����X{=�-�<�5���d~p���ٱ���	��X!���8��@ �im�O�:�����K�}�Z�k^N��;n���G����5m�W;z@����Z�e7?���[c��)�F�1�"k-a�.w�-h��5 �#U����b�T��3Rd���$�̝_vI��e���S TD��������f���R1��|�%���Xy��ǉa�H����s����� ˞B�����}dKd����1�b��Kzd.�.Gr�NVk���i%U뒺F]�H̜�6�|��,�J��D���ott�%G�4K���B/pv��t��k2�,Q�lf���\{�!�yQ�o@�X�?��f�܄�#D�~I������ŽC�Lz#���HMaA:�)��s��^\�9M)��V��i�f��=P���{�t�,����������]g�]���� �<�q��r�%4�loQ���Q�u��'�r�I�q���6W$�䯆\G�᭛M�?r�].�x��.QT��2sX��>޿�*�Ҙ��D������2F���㧕&ʹ�^_!Xh����ʎ{M�h� ��r�*`��6���6�ʼ��5�{�#'���<_��ښ$�����[�i��ax�� '�T�tI�����W���7�����=ꬋ����dO'X�Y��L��=�''t��{����T�\�b�����E�2�en?1��۷����C���O�i��^1�_����a_r��ϩ�����L��6���O$0��^Eh�����.Z���<C�iM
6�Ra�B��益3$�ޓUC�Y�&o���r?æ���-��{�`4�:Lap`ӅV�o�x�* We�cSj����E���f���x��r��~��b�/���f9d@c�l��,�j�~�e��臗����/k��8�b���瞸� {�J�t�K��g5��E'����F��O�y�62�P崛lȷk�a�?~����lہ1���+#!���\��	���=3�%�����H~k���W�N�f=Ӝ��X̫�������Å0��y��Q)���ES��=ȍ"�l����}7e3�?؛%%bz�+�G	^��p�L�6��6|i��0�}��~��������z��$v��X�	W���pj8��e��3�N׹�V��6�@���y�`�*�@�i襛���?IJ(�I!��So��b���!�	�3����������#�N<�� �.�A �{Y�Ϊ�cvz�yU�c��$����Ht��=9�b&݂�A��ǻ�g����0,[��7Po��\���܅́��/~�~�UJ�AҼ}����X����2���e�W�,�M���u��'��i����<}yߖ��An]�Ts��Yz.�����#jA8�'��s T� q��#x��t�YA������-ܰ����"y��K��¹�4���	��-� B������ߘ 
��9
��N��}=�$N��"m�����x�h%y���GFi��f�!CTh詝n�D��C�~��U�-���4��P]��6�J�[�@]�ɸ�v̻�bz�w1�6'u>�J�RH���>Y���
&L5z��!�m��t�r��eL[v5�D%ع@5��ҭ<��KB;���>楏rw<_a�в�9��l�id[��meU� ������P��٪�:{��F�\+F�?4�� �5��_ 
��"��|�AM$��9]x��-�0ku\�5Y�V�i~�\��,4���Pר;��W���#zY�Yv�s��a��i!� �GqW����1Ӑb�U�]K��b�8���8M��I�]����D����^8Q
`+��?Q��u��*9����@ F���X���>9�G�aO�*�t2$ߤ�[��C�')��H�5C�u�����/����@���jmK���}�ş�ޡm�$��iE�9��G9�Z��5����d�����z��!mX�S�܇X�`Ep[����y�$��H*T�Wt@6ݷ���Ƕ��@��?��lY���)���?��;0�t� vq�Î��9R�
&��_�㍑Թ����Y��m���P���t(m�� Ӟ>ڤ�>b��m��	x�u�nODv�9=�I!�w��+as���F�����_���w'ܴ<� �������r]���ic��yP��L>�D�:;��\��0؞O�TIԾ�F��~L3�'4%'���01�NO�����T\����:u��fn�h:c/���~�Nj�cuO���ޖ�"a��dFt4� ��ӥǔզߑ���j����hT�B���;F��������_�~�"�ot����7Ǳ��AE������ԥ���$�3��&��,��������ǰG�������2�g��M�Ŏn�����߉%t��x]��'����5Fͻׇ Z\���2����¤/�\�)M�(�|�i�!��ח����I80¬ƫ��m0_=�:WJ����A���[^u�������s�h!b�``͆�F����n���Z+_&��ol��.	�5˽/58yhM�p�}��~�Z?��%�Q���F����F��jF��:J=�\��B���� ���̝ߦ��G.�v���d��`��b�n'�W��ޜ!�R�b�tʅ;n�^���N�˅���叇I��M.ie�V���[�ʢ6i��^ �J�vV}�[���bRc��O욜WH�H���ך6��iR1����Ag'��wR��4	��P�EC&5��oC�ʚ��wa�EϮ��Ԥm/��
�ڱ���2�H�i�+5�W�� �^hxFh)5�wW��āP�,B�<4�Rљ�N���IRD��r����4Զg8�Л>���qW�(#��)�sFN�$�*]3m�R��R�k�
d7�n��,"B�Y��+�wsx�8��T�� �mr����#��l�_Q�e�(M^�zxy��#j��r�����o��#���(ۆGxu��j��u,v`�`�N�o�{p�!0� �U��>�a)�Rϗ�5c\�D�]X���Y|�i�kF�xݡb��|�[�H�9���R�)��v�����l��xjA���/��&���/Mُ��j���ӠP������y6O
���¸�H��,l?�n�[:Yk��'�Kfk�\V×b0^!��`�k��+����+{�V�QN�X\���h=ô�[��.(ӹբ��敖>�GU��ԩm�L��E� W��z��ڦT�yC||��W�!�X��fw��2���F
>  1 ,�	,y�(@`%P��`�a˅��q�M4a���8]�w��P��Ϸ���.i�%J�[~>�3<o��30��dkq�C�����y���$����b����r��h	�*�%%b��9NQ�Lu5VI�WFer�G'�\�(#�Ӏ�n�K��sb�Q����y�U���!��]wxU����e)r�qı/nx�i��T���ߞ�Qd��U�C����B�8r�!���bDû��27ƴ���=�g���Q��]���B"��&���ѠJ��3�W��J��v�$4!t#�)E̝�q<`�LNi.J&�Gw��ȕ�L:5�h�m�Iy�𤝽